PK   F�X��=Qb  �L    cirkitFile.json�[�7����@y9P�6��m�'�nl�@��c�u"K��&N��_�umuS*MՌ��d��.���[���q�(~���j��w���r2��n�����Cq�k>�Ofw���ϋ�����c�{����g����|�g����%�Ϥ��L����Ef�SM^4�d�.ݼy;~tr�K�q�.�ɇ祫TՔ�(���*++�d6׬��Ykl�8D�*�s��ZV2ϼ&��ՙ���X!�暕M�C�9kL�Q9L�%&g���!���!�Cv2��eL"�+dz�Lo���1$�ǎ�H�8�?��#��H�8�?��#�H��?�]d ��e�L|��&o�J�5j��P�aQy��9�%�.����L��d�LV��d^���Wʗ8�d���ڒ�j\��扼�`�rE�5�2Y
��d<˽�4�E
��q��W��U"gT��Q%rF��U"gT��QrFU�U!gT��O!�SH��?��O!��H�4�?��O#��H�4�?��O#��H�4�?��� �3H��?��� �3H��?��� ��H�,�?���"��H�l�?����H��+�ᜡ�D֩�t���:�� �w*g`c!�8�h0c��p'�h���Gd��Uj�~T �*E��Qc	��a5�0T�(�d��0���V��5yU�,��Ȥ�.sVI�yU�Z'	sy^h�|V�y���.���,$����J�<Eȵ��� �S���f�SN1`u%\���B�tB�*;�+��M��R��g��Dfx��(W�\��2����.e"�ez�2k\�$+E��G�����|A������+q�k(DΩ�Vvb$�#OЧ�C��)PΩI�v�
�t&j%3�~h�Ree�����U��95�Ê���)�(LV30&��K���U������R�#N``"��	������&f, �v�����'��CFX�FU9K�E���e�rDީM� ��N�x��pLި��PÊ���S�L�wjh�v��A�W��	f�fE�U��x�y\��,�t�.
�Er<N��B�\k ��^&ȼ�*3��댤'6�?A2����2j�����|:_ ��G_��?� #��I�-2jq*�E�ТZ[���{	Z�g%��b�_3�R��I�:�ॡ����h�e�F��Q�i�543�9Ŝh����P�i(�4s�9Ŝ�bNC���X�P,��4��b���k������55k�Y�4�fC�m\�Q�R����(kZ�KS:�Y��|��bSŲ��ir�j���b�)1Gw���()�ĩ8�baM3K��XҌŒf,�4c����X�h�bE3+�Ŋ�bEC���X�P�i(�4k�5Ś�bMC���X�P�i(�4�ņ�bCC�����Plh(64�Ŗ�bKC�����Pli(�g)����[C��Oo<��ڧ������oh��z��5��eB#�Oo2��Ƨ��{�^����и�ӎ	h���z���nNn0Z�z)���AC:O��<m4�2�R��e�Q̥z 4�-а�Ӷ@C���;�F�н���Ej&���>���ŝ>u�����>�4���<�@#�Ү�m����9�Ӷ����X�Ϲ��Q[���� ���ip,�i�08,�tKA#�b՘�L��B��N3�ȣ��,,׉f�F�.4"�����ٕh��\+��ԙ��բ�"#u�Z8�A�E�hQ$Z4�C�Œhq4��KC/������h f43�ÌbFC1�����4s�9Ŝ�bNC1����P�i(4��R��bAC���X�P,h(4�%Œ�bIC�$Z�P,i(�4K�%Œ�bEC���X�P�h(VD;�Ŋ�bEC���X�P�i(�4k�5Ś�?AC���X�P�i(64�ņ�bCC������h(64�-Ŗ�bKC�����Pl�R���k9�N�H�������k9[/�H�������k9[/�H�������k9[/�H���m���k9_/�H�����#u�Zhl9ۏ��:x-g'Gp�^��8R�����C@�4��?G�G�����9*<R�p�^���G�൜_�B#u�Zm�4�m��Q�nR�6��z<�0Y������|}7����_�n�����s%fe��9Qf`}%r�_0�LΩچ��� g��������m�-��l�oz&����[��� �%�������c�9�p��r����I�g�n
q������,�9�v�E�̘ѓ?E;�o�F}U[���w{�-�Ӯ��#Tމ��QB��1o1\�ӿ.�ī��|��:�Qᇘ�Q�Jr� <nAEb�F���Y����J�^�;T��۷[��¿����bV�9�#?���m�<e�s�<Z>_��o�5�t��4�9<0x���'3 �y�&��e��B�3O��N��<������� �s����t7|?� �;����9=<�s����9i�s�z�5���<P�� ��������7���So�S�ޡ<����Y��[��U���E���;�[�u��W�XO��C�U������k��V,��lw�����fs�U��aRco�Cː�92�@��Ay�̺B��%�,�����a����A��{�e/�^�ŗa�m�VQ
V��*0XX�D�%���Q,�K"ǒȱ$r,�K"ǒȱ$
,�K�@O�XERg�YX�g�Ԇ~/ϑ��u��z���6"����q}}��"�>�rM��}�E`{�ϑ}�-���Cm0�#�Ď�;RK�H-�#�Ď�
;R+�H��#��
K���$*,�
K���$j,�K�ƒ��$j,�K�ƒ��$j,�K���h�$,�K���h�$,�K���h�$Z,�K�Œh�$�$���.|S�Y�e7�u9��ز|��Qa�^�=8��_��ÁoƁm��W���|W������]��=�H]�} �FVw��t����{�pA�P��W���߹s�-u�|�H]b����|�:�<@���Z|Sϑq؏k�����/�!lفS�w�k}���>�����x���H*i`�B�7�>�c��G}��`�b����& X���:�M�o�Ђ��בu�e&�� Xa���K����z��4��L���/c�d�5�y3��X��_���ho��X�mK����A-�-�m�o)k���]�v��nuxL�c
S��<��1��)DL!Zsb
S��B�"�1E�aESȘB��-AL!c
SȘB�2�P1��)�/��B���)TL�b
S��B�:��1��)tL��z�)tL�c
S����&�01��)LLaڪ�)LLab
Sؘ��6��1����� {�~cư0��h0!d70��P�'	 k�N�r��`��I kI�N�2�v���i��a���V�0��,,��r[dUh�R�<TdX�y�H��a�<HJ�2[��תp��*º�R���Y��|�ٲ�Y0��Uu�"�o�����f~ǳ�u��!�E�����\1��~ArLAp{f̾�_�(�3���ل�"0������"SA����"��*Aa*!��ӿ��8_����g�%��6�ޭ�,�����<�=\�=��1�r5Ws���m]}?�7�5Z}7���Z}/��e[}'���[}
���T}��}U��)�Ԋ�ª���}�U��sؚ��j��}�U�8}ؚ�����
�~�����O��i��vm����~u�(�<������?�G��Hn��#�y������?2�G���n��#�y�z�ضȬ_f���~U�m}�~��m��~��m��~��m�Y��l[]�__l[)�_+l[+�_-l[-�_/|[/�_/|[/�_/|�	�~�b:�+���y����5��d�Z�a�Ov�/�)V�c�����b~���o����g�?���L���d�s0hV���Oǣ_��C��_�q���a6	�����^�^�����.}x��&�I9��������G7�Ń�z_���Z=,�si�,Y�SK`I0�~���&�Pod.��t��B����5��>h9�-�θ�"�F�eUSY�kƜu�d��%~�e��&�媘UkE�3��h��-�����}�=YTS�i�7ܚk5�V��y�t������EB^&�5��e�u��%?����Hu���>�B��;3��b��@���f���e���DE�DE�DE�DEk����a�]�`̠�b�R��+aX�W��b�&�0m����3,��oX�%v�Q��a9�V�v��Gy2պ?�6�H��#a!5+� �� m�%��&Y
�ө$,_�ԠM��*���R�A�8HW�%ܑ.1,fHLC,d� �b ]9D�]܀t)�.)!�pb�3��ab]o�"�/5Dl_j�ؾ��=�ab�b���ņ��Kۗ"�/5Dl_j�؞� �}�!b�RC������$�'6@l�q��"_)1n���/�o�����v��ů�w����hR��4�3Ucu����ta=n�d�em�R������<�$�o�~��:���׊��֕�d�Q��3�k��j��6m�� ]���RYU�I�ج��Ʉ+�gUH��]��g��Nb.L��L(-2i��
#x����ќ�Ƭ��~���*���v��ٗ�Żɴ>�̍��i�9&�����*�5ʅ)S[U(٩��b1_����C-���u���e�p>�y�du�V�x!�-/��?�&�M�@e�D��\^g��mV�B�<T�vS�o�/f����,���7�븵���ո���uq���\��%�br���|��k]/�r�y�i��إ��d���	��q���|�Y��3����0N����S�"̳�7*���2�dIaY��Z�q�a�W��y�6�)�2gk����Fj��y�0�u�y�e&�5�D��,JU繩�iª�_oG��'��ү����>��ή��򗫐�������U��z�~|��_-fW󰵽	������iM��a=��l@����b�����֖��S_�ZfZ�?���h=|�-��^��؇���Q�m���e�z�z�'��^}Įŵ�`�'���!cJ��i�ۃ���X���Ì܅���/t����݀�b[���w�
QY杊�a��E-����8Q�=�w
��N�l�SG�g.�ށs.����.�lW,�nSq���y�J)�ى��F@���Cjۀ��@Ph'@a�A�6�!�7�መ��y	[���?	#',�U��0P0�0͇	����4����h[?o	{z�~|�uƄh_M�â��rEH��
U�� Waw��|~��0�	�Qe��U>�c^g�R��24�s �@�� ��8rJ��a�*&�5s��e��pu�k�s�'/4�(��e�AE�$؀� `���PUDj�;笭{��VjO�F�O�(xb�nǟL�a�ĵ�Փ z�2����8;^��8o��0�E�e���vch����GZ<>�7� ��3Au8��q&�CP;�5����ϑ{��7?~��_E�|�㼜��!�XX�:���V��q>��x�ֿ�T��U��ɔ)��j��M�d�B����uv��7�V��ǓX��(c���Z��VG�'au��MY�s箍�9�:b�����t�R\��T�|SefmI���l<3l�r��UnwG��1�f�&�K
���E��Jaa��z�pϹ�jV�Q�l�4���vJZ�ILo�9��bc������Y#��4,A����Ub�ku��Ú�˱6<��)�M�ٵu���X̎C~����Oȵ�,�+�nӇ�z�}�Xӟ��4�a3��q�+��e�o[�}G���0Ͳ��*�y�W�xfy�m%�c5l_z�0z�Ï\�	��ɹ��\�BI�	*K���ae�^]�'�+�[�������Jn�k۲pA[W,t�me=S5�ޭ�d��)����[M�07���n����oa��z=�M���~��/:snoZ��O��d��A��v����&����ɻ�G�tr�b�.�&�?&�w�vyoNfFeQ���b�0�_̧��u�ޘc�}ѿ򾖼<]�}��E�-�P&[�]6����}����0U�?mu3��^O�������F�IM���?�����8e�Qw�2L�.L�6�7lt��ؽ�{7�4w]�
ӽ,yV�	<��2�[�iσ�R*o`C����}��:�w�P���=�)��0��������SÒ�2�rms�ᰟ��ª�'��܅%��T��_PO�q���ޞ*����ͩ����k)�ua����|:i�UÄ���=׌=IW������F�EW��(�9���U��m���q)~�0�W�
m�(����w>���k�y�ͼ�#�o�i�f��*�w��z��ԫ�_�~�i�?�#��2�m�1�;�ڀ���"��2
���o�	�z��6��Y}R캛Vբ��Ҵ��[:���0j�w��������Z���U|����כ7���ӟ���O�E��I���nG��Ƽ��gt��1/��lc­��1�6Sۘk���bB�= �sOك]f�=���`��|x*r�=�=��g��2����28Hz��l3m���0���A{p�����a7��v���/0��Xwa����c+�4;��=�����v���j��{��������;���U#e�Ö]�{�������Kۼ�N�.�_sZ��jK�=���-/��)���d^] �1lP@�M�;(Am�����h�����e�k���<�ց/jL�e���1/0�KjL���	�B�s5��=Gcj����c��=��yV2�![��rA<d�^.F�U����|���T�m,�Ƅ]��Y�Ӿ��<x��?�1a�S�Ƽ���h��`l@C�yԐ�k���6A�{Ӂa.pm�M��<�}|t��������`B��v��V&��=�*)�!U.p�]`<�r�ó��?l̬DH��%e{��RO�B~:��%�E�iT>�G�/����vj����ˇ�Q�	�H<u�%h�R�}B��Kp|.0���]�O7P�n}�i��F�#�`R�9#5�.,�ܘE4����}U�x\�q�u��p .� 0���`��\FQ�"�)W+�nĸ�nՈ���}�:���^�1aR�=Pf!;�#�����XCVq[9�I3�s3tkbA�(f`�.��R�v�(��`۷'�Q�v�z���Ԥ:����cL�8����!��mF�e��p7�����ޕ2ç׼H

�j�Z���`�b"��R�A��؇�c����^�+��Ǆ�&��iX�¡�ܨW/L��!�~9n����p��������-�%��Е�.p�_bY����K 6Go�w"$��I%�6�"u�3�xEGݞ������/�85p6������4r���kʃ<�����ɸļK��[*��GR�p��I��mg�
�b��~%���¤�;�4t1
��"!f��ě�ǝw.=���x���HJ6�q�;L��A�8
�HA1+M�3�w2	1�`���62�5��S�����L�g;�>@)�::��I�1�u��>�J�y��L����N�;�S7����L$��]�/L���~{�R)(f�I���Q�#�h&9�l#Ì�f�����ZD��ABP0���d�`P�?ԁ�����)�#��#�Ɵ�0~Q��P
�x�d:}���X�Ť�.G7��e��ɿ|��b�PL����~���o�yy�_���W�o��ZL�7Wa�>�PK   F�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   F�Xs!��}  {�  /   images/330d02b8-4530-4fd4-b6ae-26fc03cafecf.png�g\SY�>�cAQ��� *"�Q�Q�t�ё"�"B��HG�N���'�(�.%DB�HhI !�?fFt�y������0�!᜽�^�Z�j{�]������^�n�����[�%�n���-��ߘ��I��z�73�u�,/����:��n�Ⱥ��Ս|'zJM�~�K���?t_F�a�ŝ6��<�x������ޡKw�Y����֡�i��WOt��O��3uF�.�?Jh;�@>Y��_�#�5?A��ۙ䖥�R�L9ɞ�*�4�?��Y���ﾫ��o��Wm¥nL�n�k�R[�a���u?�qxS��ҝ����RR�T�"�n�����oFio���?�q�٨�S������ׯS?���Ư�[��Е?�)QAcek��h�o&��쏮yAH���;_ߙ��N7!ѹ�/�m�߻�����3�ֈB٘�<��%�j�7f }�KZ
~~,ۣ��ˋ)ybz������N� �e��A'���ˣ��.oH���f���ʞ4xd$�U�<�o�z�1���ڵwS�9a����8z���J�2���y�u�o�Pyz`� ��b��*o�G�D۳��/ep�cҘ�ܮ�%=W
��c��T��,s��;���#��S�'�4��,�)���\�jR�zK%�p+��5�'x���U��u�G�Z#����>���ԇ
^�x�6<H{��v����"�䫇�Ed��U�+'B��"�����3���O�7�65�_��E����1nZ-Z���Uލq�Nm�ě�}�̦�Q9ec\�PsV����퀴^��>l6߿ӦИG3��	�BĘ�����p�����v	��I�Q0غ���6i/Y��&��7��vJ��x\��٭2z}�v��H�?nP�[�#�-�(�'�=z��z&�l6�xh����/�� u.�d��8'��H��/��m�j{���$�E��M��w��A�7��~[���IФO�-w��$�6�^�!<�l~tyu'�i�coB~b��X1��["�c,C��ň1s��x����3�󽿵*�����G,�7]h�4��f��T� m)KA���~&��G�g���U?�����ų[�;m�|�DF��gS�dD��Ŧ<F9E�d��ݢ���J�����홈:y�U�fz4�&���ھ7T��L�1�C�����~�����K���q迪�_�����6��!�H����4+<���F���֢���7��ߪ�)�Ѫ�dSW�.��<��[ ��)�/��;D�[�Yfŏ%}�z���K��:����m��q헊;�����>P�/U�C&<d��]=�!��1wڂR����-�J��Q�r�>d��E6P:�L��^Mu~?�/�|X}�k�'��6ɑ������]��hC_�����o�	�.+ae���v"m[m����5muk���}&�n=bx�c��l�	αck�~R��'��ǇB�G�������1���R�`�_X!8��7�v>̩U�[.�8r=Uz����ȳ�(���Ll
���<�IKj�~L�{vl��|<�k��E"Vcɳߦ������Z�-.���m����k�#S2ڃj� ��ئq��9����6L`۝��/7�͞L��(�0 �R}0�|0�yX<����G��I͕�v�?�Fr�����t�H^�_qLt��{�;]v�q���1"��	N�����=���������1��ú�7;�ffE΀��`�������B�ٻ�1�D�[�kx�:#��� j�/�:/}���PR�c��t� <D`��5�H슛V4_K�������e���0�#mu����Aڼ�	E�H�a�����7������-2ծ�H�?FU�{���
+˹q�ѕ#2���~L���<�S͏����+ �q���?:``�',�:�����{{�Į8!��܏�� �iC���\���©x�//�h_�Twj|�`C����L��OD}^m�z��i+z�z�P���l
���0g���\��Pw#�x�E\> ��E���]qGd�V�=P��+��:�ds�x�䷈1;j`؏�����O/o�����׺Eॶ|t�C��i��ZB E6{�z����πsQ<�C�;��䐘�V��x�����]����g�ͅ�M�iB���=���Pƥ�C��T���B������D�=�=��I~����:���19v� �;��~tL�o��'���B��!Y�k�c�5��WZ�D��f�܇�^^���8�a����YB�b��'�"�?z�s���P!^�IRS��p�t���6�����=g�C��k �`�A���|��%K�����W�����U��*���
�_������>�'��>��"HO�8���}J)��ۗS>���d�]Pv��wl©+���qݓB��zj����:J��$��	��pwQ	�J��S��0B���w���І�-��(.uBſv���"k��=8b��IPZ��s.��m��Z��iyb[b���fޟ2�]#Ž��!�}=D��F���<%D%��Z�xڼ<B���͒�>J똵�����q�ź��e!��ʺ̘�!�o�%��h��9��l]J�������|�"�U�c�\0�D�=�z���&f�a�唖��F#u�eNY@�Mc��~$'z
i| �k�w�Na܁{�1�c���8�r�)>.޽�kcN6���ʡ�wh�_$uL`�����Ylhય��J��X&M
T�,�.�1��־v��}����^�|�B~ν���3|�]KҦ��2�G��n"a�QY��е�G��Ӱ��'D*%�^<KF`}>�]�F^� Ŷ�1��"E��p�K�Ot��A�B֙Z�������a�w����r��\���8��Z����Qd���(_7�/$ת�f�����jQ���D�2ݨ����E-������)Y^Uۙ�B��nٽ�^�Ǌ�pM�H�gG!��5����O�9j������&���·,"�ӕ�j�w��4��z��kGSez����]�X�̠3�I��l��<��W�o��s��!CQSx��Y(������rw��ˬh\E5��Wt��̓��9k0��d _��ײ-Q���xfr.2��/8�� �<����G��?���]�9f��S�-E������6�Z���/���ʶ���h F�(}D&iKpi�g��??Y+������X ����v���s�ٴP��"�ϥ��o?�`/7�l?~�oJM�=b�霤]C��Zu�c��@Wl�B�~d��Ԗ�¿��Kk����F�����h `VХ��gL븖1��:	X{$��6}"���![}��#h��LŎ��#̞�Kk0��?V�=m� ٥�����o^x��I{ǈ̆3TV�����ŏ�Tz �b�iZ)����<��#��\�]sn�/�`K���2�sq�f9��)�+,�c���F^�Q5�=e��!-�[���q2�f�����g}�Pr�)���Lj]H"�л��隶��Yl9�J�����kj��>����Gr�zGg;B?������-�{ײ�3#2S�$h��d�Y[d�<�/+��qԹ��<��Ι��T�O��ħ���ලl�~֕�6KD�}��.����H����Ԭ��w
������e���ǸÛ� ��؉�1���{��pj���{����9���>L���O�8�s�1�)�_% J�R&+�����D�M���þ=��\"+~���Q�r}�Q�v��f�L�e8��:Ǯp�뉟����f��>���c
5N��p�4u%�n(B\�}��g/@:Q�h�`�piu_g�q輡����婬�?*���gG0kx��?�����s{��_�n^�L5t��6�G�N%,ؚ'tr�Ҟ��S=b���@��1��(����F����6(Vc����Y	���F;j��Q�'/T���Dv+yA�v��}^Q�Ӹ\̓�2�)g�\������&�w�����a�1���i�l�ZKA�S�Ez}H��D�,�Hr�W�}O�E2�R�R!W�X:Sm�W^^���N�d|%?�W�S;��*;�Ayt���T�u_eI;�><7P����ɶ�E8��E�iఙ�a��I�D���<~�Į,=�$�p]�=	7�H<�G�5� /^��[Q�u!,�>~�*nљhΜ����{Ո�nz@��s������W�{���GO��H�f.�������G��P�����^j��NA��N)��X�VV4���>U�gf%g���Λ��4t8:s��?�p����c	$�9��6��5t�䰶m&i���^�����i��.��4b��z�P��
���/Hrx��l_�1�\hoEu�t���+5��yh�8ﮖOj䦠�~��ݮM���Ġ�4�8���-���ړV�QPa��L�[�tC'	#K]8�����a9�؟������ج��f�/<X�E��ZbЎ�א)P���1z��9��7"b3��~�?���~��O�)�	3����dØ|RKO顊ThU��kc��=ϊ�e7����8����Ɏ�-�N^V�2Q$�cʕ���w|؇7��*���+��.J�k"<�nDo>�=�Xf�ȟ���g�5�߫�����L��|%���}���D���]���LǓ�P��+�}c�h�ư_l2]O�� �jH�/��y���/u���`r�it,�5�=�`o��
텳x!�[KT�}L`��9�F����f��ڳ������C�/��r��F�#�e��Ļ�w�ڼW�^�'}A~�Qp�=ͩ��U��s��\�����5Qv�����,R�	�2���J�jp���8SLEk ��L��N��k:G����G;��#a;S4�j=Mlw�tﵶ"�MX�=����)�Z�u�a�E��"�`��f��ڵ�EM�#�$�S >p�����)�b�X�-l���^h����q���| �Û��v�&U��(���
�c�h�}��.��`�G�D��d�R��H�l���y��D�����"{�3g!8�YЦYH^��Z��6Jn��>��9��:6��Ά��0"��,�g�bה_om��蔞z({q�U|�\y��n(��P.��m�C�iΦ�Ѿ����$���}�v�{������9��؞T�b�01b��W��N�H�@���B�=Lݩ�����c��I������U�_w'�%7�X ʛ[+|��,SQM&t�/���/��:��>H|�YMҺZz=L�7�fU���
�_�xE�@�<�՗�Hs@�r�)O���/�rq%��*���n�o:�K�����(��W	�J@I��v�:�[*�V��󙈮%�����;��F2����Wo��$Z��B�~�ҵ��NT�h�S��}���#��(��8�dc�T�_�bئ����4A��$�Xs@�Z��/�&�����e��[)0��0��W1��D��[6�:L���s	�ӊNw�;��� ���r�^�%{�Ȃ��]f☷�/��e}�㺯�{�bR��B�J�p�n�;������U��, �ژm��1�a��ܛB��!��UU���e¸�Z�]�����粧��,HV*�$��e�y�6a&?�1�>�?�N�g.�q:�P c�ѕB�p���B�z=�6�6;r��x5"BpB���⏚��>?55�Y���K�i�aL��CK��f�l��b3�|$��D/��g���  p.�U-��.���E��e0u%T�f#�y�����3���)�V���?%�xHۦةL��t �,Qէh��6p����}���i��@�O�01��>fn��r�vCI���lرs�!���t�[7�aJELє�p[��W��u��8[� �Vy�ի�ln�}�����L�^�2����+^��Tăx�R$�r��
/Ȍ�.���� �ɵ�A5NΘ��9�Q�����Z?�ż����+_�7Z�z�=��`'Ϫ�;�Y�%�K_�yV8Z��F���̳�G:؅Ӳ�聈,��G��φ�g�M�����ox\br+�U 9i*r�-�J{�Xt�_�#��F�Ю�e�kN��,�3�{
2?�4�gIp����]~I��&莑�IK �0p�;Bi�kP��=�[E������w�b��^�~��������VS�'�}�) �_�J�t`�"�[1�9rk7�В�P%[MZZR�T��4��yL���<�Fl����k�������va�鈥*��;т�~G~.��D��u�wK�l��R�b��8�a��������\[m |�֛>o���� `!��S�j;�K���i�<�m)��T �����.��g�ʡk
�zx"�`Z��ߗ>Je�+�0�r�H��)Ma�_��2/��#��c$y��^ݟ�zc�n��8��hKó�"�FN�8���o�$�/�, S*]̨H�l'}��GO�]4rh���<�M�����K�,ܥ�=���n9Db%59�4�F���F,s1����Z��#�L�����!f�<`ʷu�����tPcR�Jg���j,����DV���#�{�B'r��0�n+���%��Ⴒp��r8$Ɠ�ĩF\�cE�-����J���ګW�ty;7��3�:f�2I`�N_�]Wz�vH�p�	j$']���>@X�Ufy���3�C���$�B�	��'zjmI3��
}�a<c�q�;�[CܻC��ͣ��]eD���l��&oUR�=������W{�64��T�ڳU���/MЖ/q�rʁ��R2��0|�h@DD�g`�����F[{�����|t���ő�
4?i�b� ���?K�F�ik2�ُV���^�'�ـ�v��[e	Ω�����O������^ L���2�5⍱�^�O�Ea�*7Q��i���v2����H�I����>�!R��a��87��1��$!�gѸ
e�-*]���q"Z	�^�	ā�1kɁ��f�y��8pi��S�aZ����q���|�fRC�k��
��I�˜@NWD�l��Fq- ���af�}g�(�؝��á�U���S gk���J	`ߌ8l�N�����{1p�n���B���e7�h �]�����Ad7=�<V��)���Mpa�}�Y���E@ �	�,�@G��J=�S.�,�~����<��4U�J#a��o��_sF>V�4l�f�^�PW7��"�R���F3Ր�(Ȣ;�sk�ҌS��7`q|g3/���������T���#)�||��}hޓ���*��� �rw"��J|��et@��aM�p	+��U̚���e�gz؏����y�1Σ�&k�+n���WP��l������y�~�VtG\��⤱6�� ��˕���a�{)fzT�_�y�£-�]���6X�r�ܭ9Ie {r�jP@_�@%[�r�?��_½h����%�yE�;o�\��S�|�F�.k$o�qd:�$����~���µ��y>�A�o��(d��(��ئ���6�୼Hc޹[7�I+��rr!�.��ҋ�˱ϸ�S	�m�(���1%u�5�W���q��Z_[Т�Ze��Aw�jir���1g?���9�B5n�l�~�X`��?
er�q�wLME__l�*�7%�b�7��)J��bl������K(�t4���o�����vq�vqX��aa�:Z�)��%�LP��a@�]���	�����hB1jq�K�X?�+#;r�b���t�-�fQ����neP~���%���L�����6O���+�Z���M����4��,H�D�D�LJ��`��V�~u��!��o
vF����*0~3�5P*�]����f�o�x����,�UZ�>=ųO��F���~b꥜^¦GwNΞl�&�8��Cf���x/|�~v�n5�㎿h�`&���'��`�t�ί�i Mej,�^..)Q@YgW�V��]�w�о���ŏ,�!��&��L������,x��� �G��0�`��(�ab���=#��6���J}c�dL\'�2i�u�!��c�L�4���.�"��':cf�u�=��ϕ��o5���Rh�o{5�"��*\���d���?U����#{.�Z�%<�4���S���㚰�~;�L,�c'�U�����Hϊ�DC��T�O���K����U�7�UM��ޠ$J����M䊗AoV:h"��U "��)�C��
�=)�i�봖����,t��o/[`��#{����\V�")�ޡ��{Ǟ��`��������~%9�x߸ޫ�ˢ�l��K폡��MpH�q���Ucԝ��S�`�z�]���k�b���di�My���e�5����+��£	��w�asw��[LP
�K�6�~���F��b
?I��r}n������B6;��J9�bEf�������u�'DVy��ug��"miT��ׁ�zX<�)^֬! �X�
���,xyV��b1���*9�l�\Sm����)7���6{��a��X��E]��Yhy�kZ��f&��
�Vz�3����*# O�뜈��]S�|v�t@#�d�1ɧ�SL��GT��ޕGQ� ^}��p�P�T�tF��UJi*�9�>�W4��GYȵ���ä��߳��-�+���fq�}|;s�Bh0	
+ǰ~�\����5⒕G�{&`M�O�����@V�@� �J8aq�q>"wc�+�>f��������/-8�)�F�Zgv�O��X�BT�0'5t�~ڸY�"�'��d�/
JS�;I��a�z6�C�fW8F���w*��t�r�a�'!U�"��}��� �4�t����X'�~��k!��P���u�ݛ�n��w�~4]����H�<>� ���r�LEl�P�79tF��>���L�!�G�)
�*f�G������k��?x�QtF���T����0Zgp�!���Z�O*gG���)yD�=_�\�(�nϺ�&�'˞�=Q9�W`#�N�z���w���qF�ܡY�R�yٗ�A���Ox��W&����_��Z��@��I�'3e㬔)���N���)�PGƜ5���i|��EU�f�2ӶZ���sVm�O�lFZĹ|]����%D�͙i�XM�wI�D�	
����F�YqV2���3~7���^�����;�y<�F�ZF�k�7�����p�e�Ȃ���������F��0�5���$�}y�>z��k��c�P��%Gl�+�&㛄�e���x��Ҁ/��;�VX07Y?w�S?jfzb��$�*�)���
�|�M+��Q�xg�S�,�c����X����>Kk��nν^����t��1��р��  ߘ6�<��#H]y����^���o�o��f���Ǟ����)��W�F�2\aK����+yJ���>�P�GF�ރ��玲�an.=Y��2�z3�{t�Hj.�\�=� �N�M3ܡ=[ �>�� �B}���3���;�2/�)2}����.ħ�Ə��f>� 61��]���>�|0#�;����F���fB|Z��D
�a����7����͡�����0m�bSZ ���ޱV	S�d����I���&E6�VH�}U`�i4|�V��8۱?�����h)]��.�s�+�����o�/&��K��by�Y�T�>ώ��h�B����ȥ��K~z�ϣ��k��p��6�� �����PAzˮ�0��N*�ȁY�ӣNiG/�]���y��yX����e�Ǝ+	�f(�*{�Ί�;[VQK�:�����N/.*����G����$Q����;�����y�<�Y(�&"9^%d��C��C0'�-:;�f�ڬ�]��;U�E4A5���6����V�)�P�pvwٓ�YC#��p;VU��S������`3NO���~�sFl��F+���N�ڲ��*��E̜g3��6��彌C/%�� �	_���0К�8f;^���,���� �H�]�z�ݮ>�җ�s�=Q��!=�A�WC�brN��D'�9�Q��ֵU�wZzJ�>c��F�B�T?�����0�����2d^r���uV��b���� �1e�k�>���hPL��_өݔ��+�%ͣ_�t�r��dy~c�P��܊���=��WE�x�l�]7��h���>\Q����v�d�x�k�`Ul���l�ә�0�t�Aͅu�v��:L�R�^\"�;O�H<�/��~ܚm��l���o#�~LF��=��6��|��\US���]�f ���ol�埰-Ev��V�6&�3p���� ^�*�I��<i��~�0�Ӆ@�մ4�S���t�tY�FƆ	i�B9j�p�]�}�{�`3:-4�ҥ�w:��FR��jP�.���(�<�J\���
�˴��J4t��gM��>���ԗF6SN��'�s=j|��r�c��V��� y�#�~*�;h�$B���a"+�F�C�9��lE�$�Ai�ǣ��@�"1]�J&=�r���J���ս�������g5`W �&%q����ץd/�ũǹ/%pZ���pI���*C�~��Osď��^n@l/Fte��a*�pl��x��fG�S���	�>%�nZ���E���Ҁ^7\�ǖ�e���=-�~i���4��!R����6I�R/!=M�r�xl�W���#�S6�6��D(���������/f�S�.���1'b-�R��}���ޔ��긖�3��$ ��z�K�JU�K$�Z�Θ��7\ZR,�Ν��C?�^�sc��&ˊ�_ɲn�U�K�G<
�;�
U_]��Dd�hY�/��<����^�~��M+kd9�ն�*��i�ͭ-+�z�E���"��so��S�9^�b{Չ!�܁�p��{����i���Bݵ�X��,��3E�V��������?
)���d��*ٟ��?��p�{���=E�	2��'fL�$j��=�)3�����6q�xWV�������Xj�vW�*"��dig�J�ς�T��fj!��ҏ!�S8�7m�n��jXZl�g���k҈��� �9���x����#�v�Lio�������(iF,��Ѝ�v����}T[�$���E��d�>/�o�DZ{Y7Y��X�R�?ۙnQ�Î�f��x5rT��Q��rw%z�6ܫ�p�Đ͋45b������*�G�em���B�;�r�`:��}��!1 ��R.��o+�&���*ؼ9��N�M}�*®��Cs��9��кw�������{m ���~̠���_�c�rwJ�FW���/�PG�ZQ֡�%�I���8�2��d�c�� �fu��e걙���D��aS���D���M��
�E�u2+����-p(�g��:�Y�^�l��gf�쨀���(��n�8�H�G�g*�����x@x 4����wW&A���R'��!��z�h��2���������&�o�#��nػ��KB�V:$]R#��P�	��j�i��V�N�",�+�e��������D��F���4�Bc*¯o��4��Jj��6SZH�R�bی|�����S�W�A<L��d�L]dH}%�I}��(�YDb��f��	���N�0!	tj���s�j�$ohUe��"�ؓ]�;Ԅ��x�x�9�����h ���Oy��W"ֺ���9�ZeL7�ۼ�%-��o# !%Ȝ�3��xUV}�����v�Z�o��x�9`C��;N.���=+J�|9���O�M�N�&-�8�r����<��2Ճs�x��,�!d������O8ɔ9�<<�,��T��:��?)<����E�T��Ɗ�))Hۯ#���}x^a9grz�C;ߥb��1bN��8ɤ}%���T�V�F._�A[~"ѿ?l��'@�o �j�0�o
SkT$s�uͽ]9�f��X!l�P@ ����Q���J86���rE?b��o��� Ŗ�_�w�T_��*�I�Rcz�_���QK�B,�:��x�A�"MqG�X��6Դ�=�(�X lRV��2����dj�y��jf1�خׂE=8b��8D|{o��/6.`
�{֪��f/U��˳tӷS���2Y�r ������pr3��D':���*C����8����)�K�0�P�\��K��Qoy��,Bw�t��b��sNf���j�:��֥��,��$�2n!]`*lTҘ�o���}k��"��D�a������FK�
_Zn7�LQ�*x6tϱ�-,�=����1uP�3{�e:��P��|��^�@���J�5�ls����ώ�,�Zz��bT�1AlfR�x�����E5�ƹ�90Ѯ�EY�-;d�k��B�sPES)-.e�P��a,jolH�3��P�3�~�+u��1�['��oR}�D�N�z<-��#Ւ��h�P�7���"�z���J9m�R}8�Xn�/ h�����wo�ݫ�eZ���W`@��[E6���0B��C׌b��PQfV�Ѡ\�%X���Mq���:�M��,�[~�jOX�w����G������t@��:W��>���Z#�U�é�H���ec��lnp,u�S��M�q�'���a`Ϲ��=��o3ǂ�i;&z�Ý���V������d<a���5�S��"KA4��`M����D<H3e%̷��G-�oؒ]B�&Y?��:(�'�fP�T�G���.�����}1�&���rX�ٖ;� �o �*�� �)Z� �]�nsɧP��젏K=���7��ӿ�
��o���D
z�.{��s��+O^�כ����x���ȿ����ڱ��A�ojQ�WN#��Y�6Ü�+օ�s��
��,����`s.E���^E�"�0�(� ��V� [%x͕�Y{"'��9������<����r ��dt�c���0��g��[v�؀Yj,jZiI�ò2B�I�����9C��n+�S�d%��9YA'c��u8���ﺒL���WU���7����߸D@����0��XHP���:�7P~s=�G�OI10�Rj$�
����T٩p�M�w��ʙ\8�aւ�[�;���Z`KU��E���H�_��P�O(s�#���pD���J�ũ��k41�欸�:��i��Z���� ��,|�j��A��)H��&��"��`E(�]�����;M���B}E8j�cWY��������4�؃o��-`6�5�M���,�^*����㶈,2]����f��:�ٮ����,�^�~��/�H!.`���o��k�U���)���E�,����z�#�{/öW�(i)��BO7g�3����#&��3NKA��Z]U�w]5��\��X���q����*9\�OE�i����Lf�<���-�!�x�V8��L��^p�;��Zg�!���ٚ���\xs����aOǡ%��3��D�D<��mp��F=;WM�6�v.������5<2���s��V��傥�
K��v�D�`r����2g����:Ǘ�c�
�&G8�\D���}U��*#�S����{7�����v��0ѕ��Fa��P�,T�ܫai�{�̨Upu̎�we@b����C%f�7��b�P�����h���G�(�J#`NR���d���[�Ĭ�eJ���'�������o�bݗ�w�.kq�@�1_��S��uM�M��3�
8��O} {5��{�J!���xg�b!��1��NK3�X^ˢ�o�˳sǭ�I)������Ơ�N�����@<��;�Q]�n�_xa����І2���W>��E�M+��r� +��3�v0��S�
r�K�E�pF#Nry�^-���i�q�=%�����!����v�7��Χ�<6�$��2 v�u��@/��SXs\v��8T�W}�m��3�+hܯ�{�?���\�89B6L�A�8W`Ҽ�*�s��MfT�^��FMÆhVý����D�"0&���vf�=�tL���l��v;�ѓ�{`��ǁ��u�~��	�v���e(z������N�!a(�"8X�Öy��el�'�F+^��z�Y��Y/�Wj�M�b�NA�8����|sY�d�Bɱ��e{�`퐵i]챏x���]ͪ^�z��k��������d�{.2kQ�����M�@ӟJ��PkkCcR�5�y��(I� Ν�Y���8.�C1)�}ei}����I��'�nuK�{k��.������/r)����,;*5 ��Y�ݍf��*^k����
/���_
��m\�q0R��aX�ߋ���*�e��g<�B���S.a6�&G�Խ�Ɉ��bV�5�����4/�L�=�B�Q+�.�(�h+S���s�=�SP�:�CȨ�|X�Q�� ��<ml����~_�1�����k��$�1a���rlI�_���+'��l���/����ˣ2�8�˜�Ղ���wpox� d{A���+C7Z��U,AN.��,���\i�]$��M������7�/�f1&��Μ&3�W�|�zCL��w|�{w��3�e=.�VIj��X�hv�p�����3�).����WXs{n�\i:��av�JAM�Dk�j' 葡���`���J��<�<<=m�U�w�N��zL���H{BI�K�}n��˴��L'=o)��/�,����C&_�VŘ~����F	�mS�I<z���+��D����[L�iby|��,�D( �w��������L��h�n�SN����j�.�R�T�[C�b��^��4��mĿ|/8���\��ޘ�x�З�z��:z$1 VJ�����ni&[,@u�>�����/����?J){>�9�e�ҺE���m��a�ki6����D���j.wf����"Ku�����XU؁�t�o�f���kJj�>�Ք���K����g;���3�9��ù�{�@�f�,��b;�ٺL}�/Oda�sG��)����I���i���Qt��Ia�̓#�5ɽ�&�l����$�e}�V��?* �B)��etfGA�^p8�^i1��,���N���7ݦRs1�)3{[��[��F�#�����uAF�@���#8'K��Vae�}K.�0�e7�\��n*�2��8��U���2Ig+=�&�\:��ɉ2���8��]F8��Yc�~�ҥ���φ}v+]��ڨ���5������ ܋���?[���o�����n.�#.o1���%[kj��.L�$}ȼ���-�r,An�@]�mX^�Z��	���-��3u��
)=�cGe��
u�N���f�;�п�4s�vu��z���}ZB�i�b��/�<��p�Iv����qh�P���u���O�D�喝۶���g�G-v���h8���I�n�fE����V�`��JC�h�P��8j�N��^ɼS��f��ř���z�%'�������C��� #d�"5"��+k�+���p��1K��S�$�m��Hiv��q �v�]�������Ķa���-I	N_�fk��h�E&�KL�ǹ$[9�ρ9_�dg���I�~�c��X�����Br�\��ѥ}t�����~u��:�\��3Fd���~�U5�#c]�������rx���s/�p�P;`�35Q����e����{�&���*o;�a
=��OyvL��Q�n���{�^�fWj5�_��Y�u�;b���������ъ��9j�Zg�*5�[vd�K�j���7�֚��`@0�#G�\�^�^�����m����ۓ�2qz�����<1�L�W�D����[h>v�Uj�7��Kv7LA*K!�0;_W��Xt8��=��:gzQt�;<�0Oխ��,���L��	���A�~cӨs�GE�%��3���Fe�l�(��������ǲl��/EV�xh�u�{�zb�yT$+M�����Ѫ�N��Pn�)��$sƓ��O�vd�
N���4��D��j�F �&�(PW�5�/�(h�tb�Ӫ���d��8:ണ�@����i�F5{��L{�@"P��N	�ꀡ��Q���9N��H���m�s��$ D�z�H�n�GP%BX�&�d��1����!q��8��<�����\c��
l{� 0�W�{��;L=0�m�Z� +��	�#�${]d��L��.ʏ7�њ�~/e�O�R�]��̞��5\���wɖ���r�y���.�e�雓�� %dpU��a>3�k"�	`y�e��p��3�Rr��#�-oD�<>0��-���?�.��#y<��X�ݾe��J��`+�⯃y���W���G�L��-!3q%ں����z��bU��X�,��[��Z���:@�JlM/���c�j�8e�WS,���vik?�&V�Ŧcf��x�C-���"�9$q%s�6����z�H��IVK�v�p����E`ڛ3S����'�'@�+sWW���ڳ���)  2އۃ��S�57|x:}/�0㱽�w���9;%P.�W�{�����Yb�>{%�@�Y�z-�r"4���1R�؁2C1Ziy֛W��P��_y�K�5W0�\���5�����E�0R��G�S~���u���{�Ym�D�~��,Mz]Vĥ��U�RZ
�\"�7`.�j1�: �\��3�>���e_RUś`��؏[J#�wS������·�$��PV�)�I�<�@��d ����������%�Ly��>�5'�rc��z5��w�����������a��`Y����+������2摠B�#=�ZңN��G���
n�[�p�pLl�"3���GҪ�\�=�z{�*A2ذ�d�/���p��^�r8��(���``C Zm/�f��߻e�ջ^W!���~���\�����Ϳ�F��۵�y�}~k��7 �<��������n�^^��_�F�g"�"([���o������#:n�<9H�y�m5G��C[�~�\��u���v���i�Xj��'u~�O;���^��>㿇���*��e�$���,�z3�yZ�Z�����TXE	����U�M��'m��Ts�~"�ȕ��ϐu=P��㾓��2��h5n�)���u!%,�9���U%Ĕ"��ZqkX�;��*ؿ�p�)ͣ��N�D:2� l������T]�	����,��~aևP��j��6�Yp�d�ٹ?6�ǵ��\4.8*��M�7�������1�'[v�fEv+�J�]%�,8������7zy�6��#2Z��y<A.�y��������J�ϭ�����A�rW����H�恵r�|/*��u��OJ��ۻ����"�Vf��	��7�k_���i�ʛ� �ڸ1�T��h~��[������!_�<K����$�lڑg���f���.�|�#��R�O��w��v�^և�Y�T��ʍ�je�2��xB��	�-n{�������W�/� +�J�s%��5�}�Ӳ$ul�}8��Į�Q�{y5 ��&��|�l�6h/�"7{�ȈY�*��d.| \�,fHZ���Z�k�e�8�����}�F%Ky{����ݰW;���5˧�Oy��ɳΖU.����~o���*�l��E9�xyKV�ʾ՛������Ym�����p�B}8�I��E��έ2y�]!����@�������	"ĝ�I���Cg��E=[��iqa҂��uvE!����r��Q�4m����i�y�0E���(��^��&h��}C������ۮ8|�B��7y�:6޷������8�o�g^���k����H�7^X=�U������Ce�����u���{��̹e����\�-z����Ko?��{hԋ���7%����BW�-i"�6���u�����{�M�%;��C�8���NgD�N��3���]��vĹ���w1�a<��!!���j؇'�0�:"5�iF�����^C�s��j-q-�Zf�fP#��6�b�<��D6���=ev�I��Z�d�����d7+��C�m~���y<�{�\�}r:D˩,1EQ�2��Ӣ$�)	Y� ��e��)[����M+�-��ӡ�`��6	31�`0��\�"u�ݿ������q�?]�1���~?����,s��BXq��}a�7�W �U۩�rŪ=�V��8޵����8>����wy^�j�w�u�u��Ā��?��Q8�7�7�9�o�3�<ʉ4��!���4��K��>@³l
JkL��nj������K���G��5�J]i,��t�i���b;`�h����Qkq�פp�Z�	oK6�̈P��>+�{�ԩ�?81�XM\�$Oǧ���p�r���� ��$|Md�����_U~F�Gm-N�8t%Z����e㡟�1�x�^��/����nY��:����/~G"b�L<)��O�e�]�<= �2�)#m�F����X��]������oN��g��\oG���w��6����-���6̾ن!��G����V����&���Y��QF��w��	[��a�ؠ�W@��7��E��܁=o�*\9�$��F�_�8~s��%)��/-1�M���sY��=�����~�1� _����K���w�]��Nߥ�вu@ٜ#���]�	軔����\�F�P��B�s3q���|-����о_���� ��^�Cl�lї˅���|��^�\�u�Xq�=Q�M�D}�K�W ��V���K_A߅�%�lUЗ8ޞoկ�c����
U���k�+�o�Wʨ�;��)-,����Wo#կ�F�u��w���~�']�.O�:��b/؃�G5?������b4ӛ�eH���qGoWN��D)׬�ެl�V9[ן�e�Gy��/��hL�)�O��X�>ew]��������k��dII+}�A�ZpMJ������<1��>�q2��-�k<�	-|�w~0>>y��ҡk��5z�M���E�1vQ�f&�u�1�veD�> q?M���27��0���2_�z��UȡI�#��]���m*]v.h��@cl��WZ�4$�� �挴*���XVը~��w/y�{�?��>5�^�{Gb�Tm�����@/ѡ���h�����=��;<_�!Pnr�.����L����C���Fn����-�Ĵ�cy���w�:{еIs�E����![2B�$jNP�t���7h�O�?��"Ϧj|�}���z+���z�Nv���Aw2�G�r䘩8
�t2�rGSu�%��z�^�q���H�fq($%gt싍�]�o����Iy0/ډ'8�M�\�3�.�N�z}��јc��{�IiY����m���UZ;�d�Z�k��H�}�I�9���r����3��NF�2�C������]�a5U�!���� �n�Ӻ/��ເ�z�)ǻ%b��V�E��!��Ul����Wz�4���9��mNۀ����づ/�+�}s�4;�n$�Χ-��ؑ�J���ʡr,��o��ZN��=��n��s��_O�]�L;���Y��g�΅�$�,��M��zx�n��MjD���XSVRI�m�x�*Q��t�,����s�=;�c��sKzx���c�Oy���9ͱw+k�ʷ�Iq����o�>��G$8�vw[�S�dj���i�����\G߅׸F��c-V��a���ĔD��,��ͱ��w�Nj{�:�y�z*��j����y��o�N�ℭ@�c+�{��$���8S<bSMO�|Hݙi��}WAʢ�oB���:���]4�����D����~X��7��.��;)���;34�T{7���ɇ�?�����W���(�)�N5=#�2��1ʟ1����w��5�I�9�n[Ny|�]��X� !t6�!��JbYM�*B��%��n�}���ܽ/�d�I�S�m��U�8~�H��S�P��F��e�X0�잓����OZF��dOPl$�xݣ1^��+?�z1Wu����6H�Ϊe�ױ�.,*Z��K�v�|4���L�$I%Y�imj�\�!�>��[9��1�|�dIѡf�dʃ���a0)m���08�V�>�33��S3�ĕE<�5U��&,"�;�vX{DP�������InR�g��K�ٿW1���/�(��FF�d�ʚE��CO�e�_3#p*��tt2s����.!R+l��b�UP�_D}^��T�	�i�fk��Tg�Y~�|W)=\� >�%�o��~n��<��I��������B���%O���+��d�N2-��{Y�d
B��M�e���]���h�EUX8�2�$��7�W��+���w0�1je�W�{�#ۃ��[4�Fy��*�`ř��H%]�u��A�����^Ad�6N���^
Ew'U��f�:��$�h�E�z�!�Yb�ES�j�`N
��B<x�{8v�rC��j[���33=]ባ\��)�QC��v�/HR�T��Jm�ma�W��`�=����Blx�]�g�J�Cb���V`��-�D��xo�J�	93�[(��R%0�Wx��
5��2�E�'Do1�K���?��5 �ٙpy�u2��y��$3����v�A��7���B���V'� �> n�=�Zjb<�?ڗ{�/�>_cWAq�M?���:S׶9��t������"�S�D�N_��~R�,X�|fft�,	�/�݁�2)�|daoI�ߑ�1�� 5kx}�A��!�l�K�#�� �U��N�A������$�#s����?�z���m�yn�� �\���	���Ī��r:X+�/��"�j&F����y�ow�U�g�G?
G�Oa��8PKt���	ƙ�����^=�u���|�v%��n��mP��}���h�c�����.��v[;��#��>�=��*Q(g5�3j,J����ىK������n���s�2_~�a8a5�ϡ�o����Puy�̫���d�ۏ��T�-ܹ��G-�ǵ:��"K��]o�&�/8E��T��O�WW
��"�C��_���x�Z�%�,!�!޲�Qn�i���=��>fR>C�,�� ��P���(��ns��u��2�q�� <Yo��PTtl�`��q�E���	lgݲٔ��  {B��R.q�GF�E�������qLZ�J�ڡ�3�k��۱q��0�f�E�@�#����BH#NG"���E��:���")��	�ai"�N�.��T���� � ��G ��VY�7�Ќ�V"M�	1�ޟ�_�|�U�{v��P,=-ݖ�+[�0~���I��0v�N�+�_�>�I��+����Bܞ�ۤ���K�Լ�m���~���D��z�3d��&$��HplI�Y}3Ϯ�N�6�`^hH�,h��)s5�7�x�Ğ�=�f������^C"�o=�l�;��Q��:��s�" ��o.ȨQ�.�%���یh1R�n�Ffxn~,j����Mdz
����J��4e
P۠�,��7yi�^�ɑv{��iy&��n�"��{?9�&������㋗��:��c�.���ne-x�D�"�B�Ǻ�s�UB�P�r��A%�ᡃF�6��d��	����;�^�S{�����M��r^���53i���L�s�RH[����O�ׄ�O�q����2hĽ��MVE�ȣ҆v��+�/����~�k1���"8)�H����1K$~~���?���!�Zm�u`��_w���"�,�M87�5���a E�
�7��6Jp�`�g���|?Q:^��aE����r���C��i���0�*�3Ŭ�e��z0fv�a *��\-m76ڧM�:�)?���\쏁�4�Zv_��Gw��9w�ֆ@������w\ߴ7�ĝ`qձ�U���� �i��?��7��� ��%=�>�q�Ք��t��X�rX��&|��g������>/^�jcʮ{*9���Gv&�O��R}@Z�{�]�m�E�Z�=�X�y}jql�J��R�@���!�f	e��U�O}�����:�%��O�h� d��r3NŶL���̟Q� r4�^�:�uO��9hu,E�hK
���!����s�%`I���� �]I��f.�|���d\p����:[�o�s��Zo/��=.��Xձ� ��t��7�%{��N�S�)��]����$z�٥$cH�@Ћ�P��`���A��Sg�]��.�Ҙ�R2�RD��3S��Yn}ei��肟�C�9K�Jٳ��̫c%��a�{��n��ؐ�ϟ��c� ��7�oH�>��{�vq�-�_�����B�sQԎ
Y����n۹�!��k<�]2k�|ui����kqRچ��)�k�o�Eb8���4]��Ǭ	R�/�
4r�5�ه8��LT�AB����A��2�A��&�����(��G�)s������_�f�����L���͸��=P���ex�o���@hh�qv︺���mV�se딹@��t��b�v�x�u��1����I ����\�U �T!2vJ	� �b��$*�OޝPIC)��#�Y�FT2�$٣1����He��v��}���1~|�����n�#�D�Ő��E���#�۰
�u����C�v���j�.�{����g�@)��!*�[�|�kK���i�ӌO��'x(�L��N� 0����vnʒ��|��X���,�Wɜ��Z�L�Sk�	���s\���}�(��*R���iC	���s�oT�궪-s#YN�K�h�ެ���na��p�{�,��v%̾2����!�ç���ચ5�K�!j��C��-�Ý֮����C��l�VN�zTO��PE�^��Hʲ��U�a�+��v
(iB%"��?�FC�!�;�-��k��a�;�FSuf�#7��EG/_���A����Q'x���s`NU�L1��`�LZ�y�^V�w_���t���o�fT�
�m�Hgi��z �K�tJN��Fyfp�7
��%��v����`������Xu��]�܋�rz�(b�[�}JY�AZ��^� �z�����,�o�di�����ODl,�?f:�CTO��!0�� >f�u�/�A�̈�Ӡ�a?6���Ҿ����hE��	)�fͿ��[z2q�-��Ƥb1L-�hN��[�xh�E��J;� �y�mF�QU���..�/C��,�{�w����-o�|�"�8�
�hۚ��  ����AϵM�}�|��z.�t�2�sd.�!L����Y^X�$�Fo&*6l��]o����7������x�Oߕ��o�.���)"�'VR}/h8��)���Z������I��<�[��e��T`���c����?˞Q��7�i�o�M��p!8VM��/0�~j����R��QA�* h@GH�9�g���ʢ�W���^*��A���#�ۛ٠�[B��z����Yڇ�(��o�g �3�6.q}�is{�����TH{�v�A��B.e_�X[��F�u�v$WQ�-I��M��c���e���ԧ$�4�����l�RF	�:��?6��Z]kF}�<�lW��̵��NX�U���ow�B4��g�23gj%C���6��]�!��'�x�l�$�l�ոv�▶���W�~;�k�`gf��٩��A�A�������R�É�)3���R[Qs����}CȨ�b��v�3�Π����:3V�j��]�Av4*�f��1�\0�_`쒓7�~������$'!j�)���z�>�&O�đ���b�Z¹/t�Rs��>9��]�<���e]���o��
�h��<a����U1}��I�m��x��������ǃ�2����o��d���m��E��ֻ���s0
_C�J*�����^+Ց�uy����ټ�cW�e�M�kj�Kk���Hk�2�L�+��w���B6�z��(��>G~)`�~��t�z���UO�.�aH��_��P&_zO��:�|����:�$��6ysH �[R�Rv`D��W��G��_�����>1��Nk��?�Mi��DT�m�C���-y���3k���6l]"=���!qV[�KR/-��)��Y�)WZ7�ϩk�"�x�A��ȡ?�p3��̠E'F5PX���mz�~�4��O��AD{���_� �mʐ����:���a��E^����L��i�}�����v�9OI-nH�׋�k��W+�܁��f�=%���e��=%�qB����V���DK�F�@������)��ݬ���M�5܀��M��v�̃v�v����L��=�n`8��t���0�-:������h���ȵc}9�bM��L�+��O�TjUpő��,�}�$�/AU���4��B6����>H�c��\���W4�W�>��z�~�^�q8��n�?-�3eqs�߉S�#�!O|7<��>�T%h4ι���zCY�#��k��O;F��>>�-I����?�e�|�^� �;��������/�{['zD9,<�s
�}�Tr�ʡ4�Xo����b�$� �Cn+��'C5�������ќz���4v�F�k��J����Ʀ��0��z�t҄k��d����-P�~�G�c���,̇�¹��)�HA� ���a�7��m^j�
6�Lǳ,*���=r�b�C��	HVc\M!Gbf7¢" ��{����[Y�� }ZB����D=�훠)����(�d���x#3�5A�*�ˀ�N�Y�jrўO��q����%[bȁQV�o2��RU�ӂbTĭZ��:կRꛘ�Z=ɛ�ό)�Uu۷p?��Tig[ �aiW7o����n�d�P�p�If�Y�6x�}�
��3��A��}2�^-�?]2�6Li���}����SL:��-c^׾�9~S��gNr�&���I}�l��ô�)��(���踵�6Z�4�H��.j�nMt՝f9��J���$w2�h������<�������;$���fٴӓ"����f=?�hG�9j�.�%sWvׂYz>���	��l[�U����0��X9���~�EC$��� j�Hku���}}1��S��۬Z��d%�E^]���Jgңz���j�f�1,�=�b���dĔuoj�MN9��L�I|���	��WC�G�ҖeL�R�t;:P�ϱ�;�PX�d�j�����3�ֲ�{5�h�7GQ��,sm�g���ݷ�mB�}�4�l �Ͷ�<�Pu�� �]M��x���|i�D-����.�C��bs�����+SB�}!G(�W�$<�������h���`�3��U��~�u�a�����6��e{t�"��ꨊ�M<|��{~�??�'=|\��VY��P�(z� a��q<0^(�"�~sA�I��p��L}����?����,�H2v�2H��]��z�u�����L��OAf��H{w�,{\��E�����E�B���ق�\�	�q3�a6-�M�o=<��!����p�	���^�<�z��@����1��hdy'�1+�ar�X�	u�zO���̬���j��!���a���s��:�V��i{һ�PR�R;MD��	��M��L��:K�M�[�&(���8�f��}����,���a;��x_;��_�&&C+�'H{�4�j�N��,FZ2Yyjf���/��p�dI�u�����^��]H*`�x��:�Ȗ��_b�e{^+>����F��O�n���ݤ�������"H7������c��s�Mhi��e}��b���RCD<�0kyo��a��PD�����s���g�}� ������ْ�b��~ ��|�I��p�8�KZ_��ۡt C�i_'�G�P!�A����>p[,24�z*u�$��ޓ�꫟��ڹ�c�]HY��%_�T�6�e���/da����qܑ�V�e�i�;�:Y<�5���΂� ���-`�=�������M�gi�����qx�5���W��Y�ϔz�;?<����㲎8]�!$�_��af+8a�T�%��1�A����=���
b4����~�<�q��Enz@���H�&^I�s!�z�^)��ؠ���,.4p���f�[G��X`q��~�@|۩q��jkykv"O�\)��{�u�Ȯ��|r��rz��@z��i�G�&��-���;)<��p�{���UZ��IFQa����\��忌1�a�y)��7� �=���\�˶�d��Ƨ���]- �?x�}ȹӻ\oHX\���+��\Wt���%?�1����2�%a����͖l5y���b��ׅ6�X6k�%5���ʺh�nY��Y���8/�lr9¨я�8���o�3�P�� �sY���fI��8	�	+N�}��
���?�v���`o��Dk)� ,�ik6��?˸����
�ٕ03��lo�)/��B��ĭL�hO�|���)��Qk4?�Z��=I��Z�����Vʒ�� w��j���~zCƉ��R��lX���%J���ؒ�5>�ަ���|�I��z�؛�2P������sa�C������o=.��mы�� �O���&�鄾��=<���o���� (w�.V'��\:9յ�2"�l�	&�\�.8�7��1��%���$������q��΄��}?�	�ϿmmU8\s�xgVٟ�5���':-�Z=���})OA؁��DvK�6�=w�����J=H�PL�T�3���Щ�SOw�,!�9�%Im����]��[�q՞7�2�Q�0�k�xS�t��)z�)�v�bKHR�"0���7��[9E��#�v,թ�?r�P;h��bz��F�hߜmS�4��¦��ܺoRWp�_���г.G {mP���u��6��J�-����z����1���%fF��+wZ���c�]}�v�Tz�M���R�����b:�*B�m]�s��D:~5���kw	�mփ�ɑ���"�5' �8�*�#� ���ayB��>�&�>�47Y��y�n|��9�,
��*���!)z��2�4FrjX6_M0���C�#�`��d�Ӎ��<��e0��#?�:��.�?,(�X��N^�t�QhYM\*���p�x$Yl�c>�u�4ְ�z
(T쿨5�c	=��W�2̔��x;�����!{SYo�Gfщ�[��P6���|�rU�i�N��z�6�����h��I�]�%&m��������y�P��Y����0�Z Kc����|x�_"�VU��R��f�|��������}\Q�O�\�qY���L�1�v�
m>�)	��h�2�JٰJ��Lu����!�M][L��.��t�LhU8��=İz��ͫ �e;I �l�ԶX°F f�����l��Az�6��8u���A�0ZF��u�Ww,�����Q�$l��~5�_��rPQ;�Xq�x�,�1��%��~F�C�0���!,�Z������ʑL֮��n�P�m�m�̩�k� dPܗ]�ko��Ӂ� �Q Z�j'���UDs��ŧ@�>.��Iv �+��lMy:�����4
�Φ���D���}�ч��+�5�*B^�+^5�HDy�rF�陋�/���Vh�.>=F�W��Z�ُ9�g��]w0WM;�i�M���_`��F�S/@<&/���$�`��vk�.�{�Xh�߾%�L����\�Th�آ��xu(jK�Ȳ����r������R�����I����Ч]�����h5������~�� 	ht��װ[��$r@�XES���b�y#�QmП;Me���#t���Y�g�b��8!	�[��M-S5֮�n.I�P^W;�<46������Z�gJ��G��̓U�dwS��RROW�컺R`
+N+�i�%A57�t�k��"��ϸ� �������xu�^���eC��n, �1I����י�Hrq��2/J�A�W�����@�y�WѩQ�{}(�o;/���;Bˑ�٬ѳ�?,�u��g!8~}�7I� x��s@w��W�%�����܊��.dU�Y@��T�ߦ/��ި�)�v(�jl%�+�
A+-��~Z� no��Q�vq�i�v(4}�d�㫯�ұ��xX�b/�FA��}wP2$~�"ĕ���x5�^��yg ����dNڀ#�jUG��pcB����K`����6(!��C e��:�<n��\�6t�M��V:>��)���Y��k�榺;d
�~z��'-����;���Z��O��A��S�T�D�&��F�X�Ҳ���֧-��
���d�����**�|u/��o	����zT��7�RQ���j�ײz}�o�y�>Х�˶��� r�&!�ɬ]Y��	�6[w�� ��?iN��ڊ���z��ͺD�� ���#G}�͗�UG����y�[��E�y�/���sߪH����2��1�l���V���Ȟ?M�<��VhNC�̝1�;������PC�US%��S�i�j��w3����� ��( ���[��J\���OFO0�3��c���`��Y/�������AC��B����S0��]�(��7KNULڿ�>�U�l?-�{nZ�g%zv;XM�����]�����(����*���o�@ƀ����?��d9/��o]�~W��LEk]��(�%�Λj�'5ib�IiO����Pg�f�h˧ddY븝ˉ�i[�Q������q����G���Fz��16���߁��
�K��Ȯk�w�9U/~w@�XXJI�Oux8��g���� �eVg��4�$pvHA�?/�����i�����4���0W@���Zj{}Vj�V����sq������уW|)�`O �l�.to����dZ^�����[W�N�pe����?{R�n�>%N�$3"�J���Ҵ�)��c��A�#&%ZbjGU�H/k���U�x�Lg9L)=|��O�E(�i����V��t��%$oV&q���P���3�0��в�m��%bY�}e,8���.��S~.�%Y,T������Ao�K�&L�C�9L�ݣd���S�|TK�%�޸�9<���7M�8f�è4Ԁ�}�;���oyX���zCL �3�~�j�]#C�;Sm�H���:|DuCI@*�^�7�m78�m�����r.���+VH��� t��-�˦����>�,��gi����g��A	E}�qj���ҩpcl"�N#�Ks���s(0���P�dm��w3����f�`�t������/,5�f��o�2;��ʘ}��FI,�(oV�d$̈MeW�*�<C�Wˠ'%*P���_����u��Zb���g�
�L�t���?�P� ���WL����m���{c�]%��-n���5]�/�(nOѨf����d�oO�?#���,Ma�cque}E���a`��픣4W�ϲػ�C;y+�]z��<���z���94�p x�b �Mc9��~>uH�-D/����|hyv�l��f /� �5�^<Λّǿ�����F����x8�Z*|�E�!���"j2;���s����������~�ku������lHN.��0�{���4����)Y��C�!����9Ⱥ �`#t�/B�"��U3O,��]�ɰ�x!� vGkʕ���އ�שHǔo@Ke�ga���a'~*��Ě������7�#؇��'u/��W�:2�=������ă_<u(��c�>��'ypf�"$o������i���`!�_�{8ۚ�ԗ�v��dE�
�Y�@m+u�m����ͼi�����nm":d�Uz?s�e���Թt0�ҘD)�F�u3�#�4���[���\,�c�u�X�H��P*��`�����WƄ�w�6��n��,�7aY����tf�)}@xt���e
~_<�n�>u����{�~��BnyY=F[�f�[�=1OQёl49Qr�q����G�0J��Q�}�~z��`_{!/�ă*����47 u@�g��֠��؈�D�S��BcV���@W���剟 �}=��U�{�*�,A�V;�ց������+���O�]t�F�pFL�d:� �5uc w��&$�< ]Y/A�H@t�[
\}��B������h�~�=�1H=��Q/���V6���9�6Զ#�D5���z�ű�:VZw�R�Z������s1��.z"7UWa��F��)Cn���E���ϔ�Hp�j ���q:b���E~�?an��������8�LGB/M񧏺��ܦ��M�����ol�O.��cRR#����گ���)̤�,�tS1���W�u6��� ��]��&R�z���_�~�����)���)w�.����̴c�*j4V�g
�� �����f��Om�6g��E�,;�O�Z���� X��[^��7R���. �*�t_�c�#9Z���ԧ0p���+6���)��N�H�s ���c!A�O���~jM�BDά��r�	x���Qv�U�뭰�U���ڨ�A2�㫮lo�P�s7�g�Th����Xj|���Mh# -�"�?'��󍪾v�v�}k
~��~�懶�^F|���xYz2XC�!��o��u4�� ��o��u��u��|p���\�f���Z�~z|$����{�?�?p��"6k>X�����?>�ӺK���a����p?�~h�?\+>"�P�R�K�.U�y}���_����V�D����������,��h?J~E~(��s��շ��\+*��z��֏�$�L6>P1U�}��K}Z����w�
^�lJ_�����S�K2� ��e����Ty���|킩�L�9f��q�a�vi#z��*4�Q�����i���e���5��C?�-`�$��gL����A���w���q��p��Nl�P8#���;n����B	~wX�Pfm)�G<���6�Lx�E0���D�-��)��j�b/���UZY͞:/�������6^�XFCAz��&�Om��ε����D�aY�2����K΂�c^��=�I��{���K>�v��-.l\V@�bS��-��@���I���/m�?�.w
	 ��)�J�������$���8�/'�hsʪ���Vk�ƮCW]5��� ���ھx����X�-궉���}�K
�g�RSkܯ�M�$�5�r��Aa��1Z��/�
,�w� ���K��5�����_5�����9o&��LK=�g_�i��X�ᒶ��ӇQ�D�Mx��ޜ��-�^Ѯ�{�[��:�+c�U|�l�?]��?Up9Gm�����y�i�)�0N*���e6�cX�}G��7dF0�%�g-��ñ�vh	���>�\�׿������lv𻜖�!v~�*�S���\8$�T�0�����ս�Sm[E#sE:��N��&���u���m��{*I^o�ק��V�]|�tĞ�����5�7.�
��
DP�sG��R(&�<L�}p��&:�4���Dܮees��ݳ�"!���D�-������DR�{{��} �E'��R`�r^YT���V�l�Y`4�܅��a
?D�ȡ����l}O��)�����U�`�Mw����^_��B#l+4��u#Df�F����(��6�	v������\ԇ���p ����i�m7��sxXqʹ��{Dw����j�/�^�<L��j)e���Z��^i[�w ��uF����X��|��kZ>�.� ��i�Zx�߶A�} �� ��D���[I���xZ��u�V,V���@JI�^����=�y���O��� ;j�J��YS.:�->���@U,V�w���5g_C��Co��Q��4�װ��$߬Į�ٌ�G����b�،���6L7I;pD�Ξ�Se���/�z�`�l�l)�&қCmO2Ej ����l ���rњ����2߫q��/A��f�b�U^�a�>���|���z>�7�qr�TLm7�N]҄�@/�y�2\E?�'���I��v׷A+�$�M`�������*��]����@}l���/����l�j*��8N���b��^���0�p)k�sY
��ο�{����Y��zq���_�|q�h�Z��ϰ	}��l�?߳'��;��_�_�-�u�]ge�|����8[s�/� �3<b��s���PK   F�X����(w  +�  /   images/42266fcd-641e-4cfa-a619-b442e1b7bf10.png�|wPSo�.,�X�( �KT����t�C(�;(�Ho��;�)���Mi���йI�}�9ws�Ν��a�	�d�k�{�g=�Zk�PMu�kT�Tה^>ע��(HAqf����贂��/�߽�s��0T �;s��39
��)��r@ϴթ��@�c��~^�Sy�m�?H�����@����&%`������;��Ɩ����*.#9οdC6��񕭖Ĉ�P��?Y³�T��^Ե�y���ݑb�ћ���������.{�?ާ��<��7o$�'������������g���+S�*�%+���9v�G���4t,�
�I�@A8=(��#�2ڑ���,�����u-��k�E�Cps%�%]-
ϐ��G]����[�?ffL��#"�yd����gP�==���U�c��\�}�?u�IN�OIIy����2�\̗�GOWW�����k;�-�YϤm4b����}��Y*��h�+�e��/�tP�i.Ӕ�����#�϶H�N"�ii�H=�).�%Z����\��� ӿ�F���N���/� t����Z��N_�~���ӝ�hY�4<<:w��Gxx8D�J����ML����#O��	A��ҥXm��k+���|�*�[c1s�Qf�C	���e����~s��oZ�/	�ǥ��{����������rw�b�0�C�t#>#�����p�1��|1�8��;����Y��h]�/��2����$�i̍=��3$�{����7�����ܩݖ�%��}W<2��ɔ��І������q-ԕ�k����[-����5(���Μ���h)� �7H榤 ._�m*�T9!)���l5Fl��gR���

�_#�tw�}�Y��>=:�9��)�_O����`m�q�vM��R��S�t�8���������*g2N=�-ʔ˲↩�ު7��ˊk�g���\�j��W�7,%����L��ض��h��	�m��V���O�����_�،����^�,�7�uKK���Ʌo�pq���Ù�� �5=4�����jɩDs�!�Yݜ�Y���b���nx�����s�g[o�3�6
����?��g���;wq[�X�|�.a�Kn����{�>p����z����� ԧk�Jo4c���;���P&÷W��\`⾻a�[�)��b����FFӃN����?���Ó@TA�����]��!��%����v��^�����K�j<��/e���nSI��{��T�o��x�{�:u��7��_vb��,":��5���,v��VKN�ê������xZ~��s^{�z9U5)de/�	bQ���UmB�Tc��H����Y���{�Ԯ����,7����;�c�����:a�i�R��I�2�^�2Jq���)++K�P�ـA�MIv9U�@����E��#�6]��8��GHڝ�X��t�1�A�ڏhy۱�7�!��8�|�jiG��:_)�t��o55i5��� �*����G����cXO��[�W�_���+?nph���k핻:i��p���5dɆz��W�@qX�����|�c묋]��S3���Ɇ�4�W�<�����kj�nrg�}�h����_t�N�D�=�[15�Ҭi���cm�^��v5*ύXe����U�u���)���)�lPCP������Cz�w;W��d�/:��+۾O{�����5Y@r�,l��פ��7jK(^0��'�^wm�k��r�������_^F�z�R����1�`@�{��^��ט�����ǻ� V4}��K�6�����cSͬp@:E׆Q�Z9N80~�P�NO�����V�� ��;~���#<	��e@ɮ� =���zo�W��L�SE�2"j_;��g,�m�+��i��grg>2�ޣ�dF��1��O]�l���&^�H ڨ�S/E=|He�/"�}�X�"kTލ#�R����l�:,c�
/��"M����٤Y:s�I6?����!P�#�9���ˢ�tE�Z���cu�ZV�L����'u�f�R��״�el�y�}x��?������"����c�MjMgϳ]sHL��=ҪaNO�
7& ??n��`@��F��F���r����W�{6�G"�8�snSѾH�f��1��4�a��#�'�0�u����/�.::�Z��R��6�
g��=!s|5���t{��2��R>���M�VZ����>�� �M<���=d!�b���ʐ}�����Q�4�_W~(-m�	�C/=�}U,����u�����=����Ҩ8'
oz83�y�z����H@�ˢ/��;�ALɩ|}��n��y�wꍑ�xj8�[���u�H�{��;��7���ԡq(��]v���X��ʺ�c��٦�B�^.ݸ��o��dO,��Ua٩�2���}br�3B ���&D�h���������G&�=^Z�@�C�[�o>&u�g�:V�9�m|���Ewt��Q��҅�b@�m-�6��l����}���&$�p��=�zq�<�:w��+ ��������[��'٥�+BZ%����h����i?
�>��ɷʮN
S�`Я� 1ܿ�� ����cޢ克�=AS�d�"qz��3�h���͹����̷M�,���_�<^%L{��"��l�A�/,v�,��_���M�8�"�f�2m�V6:���*�����3�))Qz�{�`��%�!�A�;D���G��c�w.�{�9���csz�7�.W��Y���;��B��`��zMp*�H�;F������t�?�s,�C���-e�z�A++-P�3����7XĪ���~�l�F��g\}���"���î��Q�l�Ԙ�T�kǇW�h^�����y%��13>bZ������C@oݼ5�$�cr��ks3{�Փ(��Z��dֹ�]Ѽ7�������Qe@���:�� ��/n+���	�����jXD]vxU�^�&�00>�ѹj?��۱�n����"7�l^ٙ�-�� "����+G�ϩ$|q������%-�e�� r��6#�U\�����m�F)G�e�*۵��*�u�Tc��#Ϻk�Ӵ��&^�E�g/��I��-F)1�z�����ί���c�|���vl@�]񍹢���1��a�e\����i�F`՛%�R.Փ��DȞUo���R�k�e����v��I�e�7��:��C�=D���{�f|yV��TM��.��E+���<m�P�)I\G���aoh�K�������L�U�n��/��Z�|U�&�[C��&�C�8��yǠ�t��H�
I���WSfn<�)�^�v�?�e�6�ļ��ã#���-|��D�1�I�3E�y�����D�NI+O.e;6U浺n�/ ck��S�XEt� �Ҽ��Xla�cf#@̾%N"Qע�MR7��^~�Qa����1���c�ny��TM��`lTZO����z��f���G�jȈm�,j��Y�)<e!ȵ��:���jDt{�e95K(���Q��z|��N�\T #�#�פ�q��s�޿ٸ�����Q(��߭�ފ�k_���=}�k�l���JҎ��M�U�D@��r��c��nk����2&���o˽o��K���<��4�ٳ��� /Х���߷e@�0�"�2���4�<@�G�� ��ؓ�0���Uȣ���v�EǨ.a��~�-]-D��`�fAL8�������aUr^s�B���R�a1?vv��3;6���x"�P�]�o{��풴�%78v�En�(]�8�y|�l�FP	�nfE�ǡ&ʵ}2N.�C���M�&���N$
z��
wq^0u=$�-�*l6	�n�lj<�o\��]�������c��&<j0��c,A�a��p�cٓR���#@M������up�7�f��@U��,J�|��I&L�W�S#3��ha�~��p�|��H1�2��݊��OivV4�`�D)g��8#��w�����}  �V� ���T�ݑr��F0}�������p�eW���=�: *�QK^�.ϖ��l6�G���(f�g
i���#�U���uNq��
ڱ{�Ƚ�ЃW^PG�D"T+�s���������2pD3��@��c͋l�]���b��T*�����߻��.�2#���"MRO^�4�o��hQҘ��";�x��͛j<C�,-m��0����m�+��9{���-֍����4%�Ia���J���Ƭ��,[���_f�lG��D�n%pYC|���>3Yg<9�Ey->CgO����|$�7����R��B:����ˋ���l���D��aV֗�Lf���?�����hd��@G��}o���������|k.��Z�����Dd�a����1< ���#���[:^�]5��h
ɨ�"V�����#��h�ɶ�AFTl_��«HQl�}�i;��o�m��j��b�N�z���Ѧ���t�2]�ĥ��r#x�J�H��*�V�.�EŉJo��߯,�����
�O���~�:h�ie���+�Q�1�Q�O��W��x��>Q��Y�����+�t����h�n��כB���k���M��(`1�n��P|�z�P��4=��H�}����)�	N����0#�8ݫބeob;YSܪ�q�JZ�}�o�⫔2�z���-����K�
wﰆ��	(�Vy)1�b����j?��E�h�V�q�����b�^,6�[XtVĈn���]��/O�#W~��:&�'��Q��J�(��qI����������1�µ|�e,��B�,g��lQ����6X�~�r�:!o۵��]��Q�o���@s@~��jC��V�l���̛�g6���v��LO�n�9F�y����c-���k �R��ŀ���b���ٴ��'��˶��3������������6f�2氿h�7Q5�ÊMbY���]�3�����Z��Q&�O��K�-��<�=!�BӁ m}ؚ]�l�r�\Ṛc:���
�D}N���U�>�<Z=���Ũ\��o�0�t 
@n�o���l����X����w�,����
�CӿPqs����$�Y�"�r��m4�G�r�����~=��ب~8�n��DU�x���/2j�<6�Y�	�GG��H�f�|�\��̇��ՠ���0Ҽ�.6�m!�����l�^m�$��}�Ww�9h���a��J��@�$���뼴��l�C�J����d/��e�>3?^) x���M��%52k.��t�\����t���kS���W ��F��2���DpR��T��'�d�p�f���� �e���a�g�O�յ�*�y���*i�w �^�(!k���x�TQ˚��$�}�8�]�L���L�+�GN!�RR`�����pۯ�5��qOn�Ϟ!F���b��>7��i���xShl0~В��D�Ȫ"���iR���;���15"�þ�(�u��*F+7�#H��:��CI����eF>ܺ�Q��e2T:XJ㿪Ljy.D�h��ujyW���kϛz��DX��Wo@�Lϝ)\x�{z,�U�B�VV�Ȗ!��`)�0C����9��ii( ++������uƙ��t�Qȃ�_��I;�Qna��\H��/���A�O{�9aX��9��(>�F>~|9U��`���Pv��7fs�'�2�7���.2TW�s>��D���d&�	�U�+d�o�{�(F�p��&9�1z��G#�cuĽ�%Es�OJ�E	o *٠F�۽�5a����r°M�h�}6A�P	`ץO�,�������(��m�Bxc]'m���W ���!���݃=�wD���U���Rm.�U"�5�_����WꇷP�g���[�<�Y��	�jg��i��Jtn�t�,��#%TO�h�
��h�˗��H-����`�_�L>�a6��rR!ő�6��|�����d������
R�tC骗#/H,떾Y	��Yב�Y��k_B��U����ի�)>>]�
T�X�@n�G
V<�t�!1��E��1:�?
��H�W��/W�z��%�/��&.&eyW�%(�!��)с#������f�
J�-) �8���Q�S�E.*2{`ݘz�"Ea�{x�bQy�h��J�os�q�(U�4��|�X���1��&c�U|���V��f�p����kJ'�ۻ��������>��܌�n{M4�B-|,��������Ђ���*�_}R�N��wG��C�b�E��A�?��m.�(�:/�X#
�c��I��B'���+����cb���&1�%=���n����kt����.Uf�uT&ڑ�c9�i�Y�]�7����������p�;,�C��:���* ��m�a4���� h?�s�.9 [�j	ix�v�k�Te�y൷���mU��S�L�8^�,�VS��Y��ky!sا~��}ڨCߢ��5@����#����f��hj�1��������O1l���蠓��L z��ge�����Ή�Is���~�bp߱��|A�Ll�՜nk�י[���:��z�㥶#����B���'�ʨ.m�`!%�M\����a��W�<��:��rH({A����Bv�1(k��vo�GI�I�,��U/�U ���#���ILl����&YE+{�|
'�ᰱ����2�Z�?�I���/�j	o"�f�[;n�|���Oײ:���4���kX�Tt'��B�BǵTs�` י�I��r�u�W��X֦�J�ݖ�T��$=�T�,{���a�WT���5�'O��J�������\M_iY�9�}|���G�9=��M�\���hw�p��������զ�	B��4_�5��� ���N#r��'UoS�RP�b����!��cs/���m���T���G���zz����[�}�&g�v��c�P��Gc�e�C�y� 7e�t�<���!� ?~��5�q�>�zF���{P������h5ns�0��h�I@��ߝ��p�g  e�7��~[�U�,������F��#���j��0����ְp�2ouD:1p�o+�i�3zܰ�Bc�G�h��e+*�f$!_��Gv@��ъ����"�Y�:�O��﨨��|����3#�c���Q��{�Zll,�fny�	|Ks�	����+��&1�e�j���J=V����;�,F_�FLnBQ�"�{o_wԻ�y!���-)S��s1�|��39IMy`�n��G�$]IyT_w��Y���Ⱥ��H�hi%�7\�5�������i�u1��-+�,��Mx�1��`y<��*q�M����3#w���6�Bk�zm��A3��V�ۚ��-��Nn��W��|/�)9�Z�����C-�] :E�b0���S�Htq�G�ʽ�Ws��yTB=��J�Z�� �<D|�o�Wqp�Q�wo�Ņw�Fvk��BO$� �珎y��ER>��z��^n��=`6�W�\gU�ufZV��˅��g}�ɖ����W�����c�����isv����fdqQ� U�J��V�����t����ƫ
4Gp��Hy7�G��!��zX���0�Y�e��ڬ�	�̭&]�h�^wo��ʳAAy>�Y\�D��ڧ��=�?�6d�5�?s�E��&c!��F�u����ʝfա����{S�W�i�c�K��]�������j���kG�5�B�S�\}B�~���(�Ư:�[����%%��������6�5W��.]���5���먥��׮�W�����]�P�R�j��t�]��V�|Y8Zjx�~�F�x��A�?��F.�}s�o�5���<��⡫��K{���Q����f2�dO��f�O��)�M���X�Vs$7��|���QN% �)��d�@;����i�1c��2tD�6G��ԏ��s�z�j�ݺ�Ҿ\�y���(��Ħ�"�:Q�Q���3�^1��gy�^�vu8����E���?�%�Q ��D�29(�*��o���f��yJɣ�B���o�~���RT��0H_8���=n#F�NN0%��
D�x�ey�~���e%�V�T��;����tk�2����-��i��IhǣT5�7ۘ ���8Ul�4��؍-�é#8��Z㚄x���<.��C�S,�	�Y�[�r���X�W��I�9^�7 2�v�=�j�oθ\��w �s���򄋠z���$���`S���hIZ��}&�����'�i:�	_;�p�p�o��~�wQW R��}�[{���?��1��2B��Oq�&���PIk���ٛ� h+�9Yp��]m��{byΑJ��O1�c��ʼ�� ��w�VF��Ei�&��{�#���4�Qq�"uO�x*􅍾NG.�\��<��IR������*}_U��  �f���=/�N|�lF<3���O�Z,����s|���q���`nC��`EoU���C���I����P5X�/��K��6h��nhn�_�f����H}�ciO�����aCe���aM	E�Hk���l-	����"�ᾡ�-t�O�fc��Bc?�Y1�s���9����V����)T^b� �UVd�pS�o���ߘ��%����ZT�����qF>����6������-הS$�NIrق4�q�5��D^�6��B�R+��/��G���	�}u���r���X�P���V�C�� K��È�x'5.�KN]�F��_o���C�ɪ�<��SgڃT�X�&bY�n� /?�>�97�d>�ڶ9s�䌗/O3��&74�K�J��'�q uf�6�CO�I&NF��o�3d_/��E"��wxde��t'^�T�nD��&�^����|}���åo��W��_��1���Mf�z�y���ըX���$7E��������%^�i����I2C�>��04�2V���wa;� A$'#pA�1�%�n�%cz���...�t��<����x\���1�5/8vr���E�92>�t���.��y�~�{�,��)LO`�����JLT�ZKH�㱾�<v���!�J܀a��(x3w%��kz �ziZ��Z�u��s�B�JC��z��_bq]�3��=�5!$�(�;��#tx�z�n�q�D5�ʝ�J�#����>�/l��������$-kT�L�@Ña���)LhAQ��=x������|S�x�ɖ�%��)?~���{��A����T-�m�Y#y���$ӗk���ǍwD�8�Ŧ�	�	�j����<<�+�RV�&�ȒZ|�}z�fů��N��fa#��i�o�o��xab��z<ӌӹ|���W.z��l���Uq���к�!M0����	tyC�v���ZL�yo']�]?����2.�|�R��&7�V�����"�q=;�K������zy[˂��o����|�G��yǇ@r�1	���1�)�5��9
�� J��?��T���v�9�$�mNw����l�+Ýֻ��p"�)����0>��Q����a��qL��/��g(���y*H�(6��0d�>5
B��?�
u}%���i�a{���{0O��X�t$�R�P�|��;�m����ڕILO���Ui?}��H�tR��\�B�,Vc�+m0 �f�}���~�"c�&�M��a�\��8��t���\��.v�ޖ�Tvq'�ơ
n��8zv�w� t@;6�cO�p:v�l.�A�̼ݫ�|2�VL|�[Q��ή�<"�@�����P=�s�V�"�)����b֭���s-��:i	�2��.e�|��E��"W��̂i֯�׾��hy&��/�	h�2�U�>�X���d�z����a����XR���֘�,���;^���\��m!�WF���ޘ	�
���%q%�0r��tGm�
�V
�en8ޞ������o�J49�M���=�����-rl��k�U���<�	w:V8O�/�:ױKtq){��B.��_h	�s��܌�;^>�H�XM�	�o��IHS�)�4�M�'ϋ�U�{۳���ȃ	���'��, �=Ó���_�ZѺ�r�@R*:�"��K����Z����pX�ŏ�Z����؋�D��ߦ��2�ΔM�AьdC��m�]�vVl`�YMNw�I��z��P����dE0�}\��[��~>�Yz���$�ůӞ��{"<�ə)Ӆ�K��#~����^"DF�����7�+h��2�뭻�,k��wƟ��
����5�ϔ*�*���s�"�Z���X��l�ӑ�so�"PCv#�3�D����s�d�Ulr]���㿤)�7��N6�%YYOߜSIYvcv*V~(i�}��h��6~L9�M>q��9��b��G��4�>����3�)7��m���a�e��=^S�G������ix�qL=h�L�wN�8 y���i���e�
<�K-��K�lpn� ƯQHR���ML��8E|b�*a7�{݇�Gc)Q�	�ņ����$Q�9�09\ ٵZ\x}Cj�z�.6����ؤ>S��:|1f�����k���3*&��I��	�8}���7��ٰxSs�2�2���C�L��H�wwףb���0+#�Z�ۧ9a��+Z����o"��5�5*�"b������f=�B���~�F|{����UaF��[�)Ά����6�Ձ^��?�Y�?�oܖ��W�2��M~F��ZZ��a�e��ɝ%U�Id�x���~�"z�A��<�I�S��3mi?QFcNZ��E;2P��Y���j��JC�����f�)V!�O�Y����Xy�������N�i���$/}ל���l����7�댩���][�1!�y����Sߪ �03nlҜ1�6���09�V�L
xX��o�=�{\�����ڈd���s=r2d ;��q�Q$�y\n,�GS1�����S�F}�(�l�qT�ʗ����Q ��2�Z+��y�`MH	n�"ۙ�`K�O/�����8o���\�����S�V�/��{�U����.r�T�	9&�5�D�¯�݊'��[�D��
���j��>�IHX!���lS����5��L�8X��c�B�F���6���
��9wJ��=$ZDFX� 2�:����!�sW�m�9�o3>"���o�=���	�	Rm�5�Bu���"V!�G�ˬڡQa�T�B.���l�Ge�aɬC�P0��XF�o�ҩ�۫��q��L�۠�r�-��wQv�;�2���s(U���)��� A�y5�����p3�5Lڛ��\�~�c-mTB$�Z_@���p���p�����}�-������|F�jG���%�"�%���>��췦
�Z�g�=P^�LFu6j�Q��r���)��/� �3��U��G��XR_(���B.��ٕ��$2����<U��V��j��	ҭР�N�kl��}��5JF����ųU���0U&	�u��TǀQW��Ӥ8�=�d��Fנ�����ki	�mM��*AZ{�)�������e�r�LC��������Nny���	=����ņ��4_���Z]���dZ�����따ߖ+׋Y����PQU����<H-�+Ź�ǰ��ɻ�o�Z���ex[����������֪2��5 �/��SV�����{Ǒ*���)��pSJ"�xZ�٦<��6}�}�w�^
u�c�O���a��:>]fn�����A.ۨĦ�Q���ve"�םS���J�T����N2��dʹo�r ����5�b�I��	cT�!5�����3%UV����s�i\�\��:$�4�=iP1L����ã3,cEĲ1#"�ɳ����j�쥢�q�Q�}	�v,0���X�F��+������â�����@O�f���k�Q�2M�h&7]_� �O�k!Lq^���ĥzM�t� �����O�~0�Iʹ�ג\!����;>3C�A�Р�$r>�_'���U=���4����*��AU'o\�\)�`>�v8�U'�C{�=I�M˶�k�i��?��x!�O��F��,���Ϗ���L�&�����➢�9jUj��D!n�{�#��)?�;���rΗ��}���[q�*_n4��E�ˡ����{�����OTo ]�Tw<EK������!��I�Ï���U��w�E&`����U��/@�Nï.��n����5��!�&H����t{㑼�osX~k�c���9r�#���TF=L�A���O]�5����*�/Q��7ʈYŇܯp��0�B�����_�s�^k�J�+��%��w�tEʄG��=���+;�r�	l���F`������ve�Ʈ����{���梚=�-�r)�RLO6��2�?w�Cdh��e�-M���[�N�  �͵�P7��5*j����P�����<|w��."�T�?!�
��[�KBnB>��N3�"�D���(��_�S��~��y��8<�Պ�?���!�h"X1z�; ���f�\�TuEX=Ó5pzuGw!�N�$��]ɤZ����0��'km�!��Bm���O ���L��� 鎺���.��x-�u��%4忹(
C�.L�P��5�hJʓ��� ���a�F�Dݦ����!���,��:��_��v1��+���,_H��%��-�{#/�����I1:=���[�N������T����jkx�}�a����" k�r�u���/��/�"�G\���L7.���\O���
{���R3�jE6쳶}���S�c_�c�6��L$Iח�C�ܮU/�j&�x]qk�SH#6Rp��`��x&<�,���AN�I&���MM��V#Ҁ��v姱^����ɲ��
e�_�h�A�,`���b1���A��k��,���4��{�5� �	+ߞ��v�=ĜkhepY�>���^�ا�G0�P���/ז&���?�qŜL�0T�B�7�iv�9��k�����6��߾rח�:*\�,�,��
jh�xݦ�����9 ���d��Ŀ�H����Y�耓x2�&�ʅa�mKn�L��ϗrA�Qb�}5����ߦJ�r������8�W���U�w�ϯO�4��$��=���{�u�
hF.�ɜ��_�U�L�Z,2��g0�Oא�ڈ��tE�p��ڈ�����*|Ο�jS�םS(�����A;$[<��_ s���i��^���05*wl>�u��Ĕ�<����n�,����@�lb6n/E���ma'�m ���`�u�飽D�����kk�I�:����V1K�(�c�
�RH="�d���1��M�����Ot���]�⣵��Q}��I�=���-�lפZ_�0)��Sc����8���Iv6gG�G\v[�3���� �Tq>���x���c��Eg����7�U�dPҼ�'2>e�I��Ti�=��j��?O�"�H�OK��p(t����iD��D���΂N8�C����/{α�Po;
Yv�[eķ�a��������Bk�� !��0h �����sx��m�0�0c�y�c�fO���|�0�]�)>ZJtW?1�؟-O��wux<ҟ#���&E��P~��.?��2�Y.�U(yc�\.�����R<5�Σ������Q���s��xD_�0�T���Ym`�OE������fuy���}L��WF!���vN�q^��U�ׁ��%�$s��>xj��18��2� &��h�u�	����ohk���:l7ЯE(��̒�l�L�c��n����	T����'�������dS0s�Q�B@nr��s
�Ew��05�,�v���Gt2os스FИ�� K\���`kC��b�eP)+S��"�Hҝ'ͫS�Ȏ�<�%�h�y�Qn�ާ2��C�:�A�q�R�~��L�ƭ�4�<2���l׳�'���_A��2��XL�ɲ/�h�?U4uze�f�˶��6��v�q�y�<�r��q��ј@Bu2����_+���3ʤ���g䌳���t�Wj�|���&N83S����އ��DJ�W�sJG��\,��U���o�")�@2�~yU�K���ޑ�g $>��q�q8M/��d#q�u^c2�kS�3xX���"0h�(���343�(��J��
Wmܢ^zc��|�]�b�)Կ�+��%D�f��D�;�(����jY*��gm�,�[�U���m7�6|5��<]�5�]�ȷ}�������~�െ]JX���ր.:��f5o�F\�f�&�m,U^����f�gGނ�n<N��"5��R��D�W��19���U�#f�h�,.^!l	�p�Y*��Q~���S��X��4g�\���&x~7��o�ᵨ5��QcHuO���w_O@/���Y��� 9~szL�"ߞ#��L�~}��#c~L�X�/eז%2b�&w�&yM��7^��̘s��/{[:gE�io�O�#k$Zb��:Z<��}��	-�r�U�z�ח�|w�����p0�V^�IL=�rJ����?��ͱ��]g�I���&��%$���D���@��Z��fK�|�)	��a��`�O�0�`�t\�CGs�q$�����x����-=�m�}-}qY�~�^G�=Z�Z�]q�<.J	�j$"��\-?H� 2L`���p�����'ہ�=w���
@%�*�G��0���y�³�$ΰq�ּm���wB�����כ��醩M�_ۙ�=QG��� 0�lP�@�%�m>s�u���'��<� M(�?{n~6ߵ.�]��0_���aT�҇�_-R�ɾ�Fλ��l?�¨Fd^�;�uTZ'=��,����E�S����1<�o�D�������F7X�N�	k%kuz�!�^W�=�P�S��ϗO��(�2��� {}Y3:s�M����8��q��*��/��y�>�f����y�)��2��|yvq�)kJ?>��
���˹�ʿ-N=��餋|n7ļkH��u(�V(�{�α�.2�a�ٳ��Tf)ǽc ���ǖ�G�RdD��n}���^��{R鱧/@9�5�-x��[ A�4���(hC�Cb��D�<1�Gmɐ���)�T�����5*!�rci�������m���**�9�E����b���0B��n關��z7�Q��*KY��i'�s�]��!
#S�v��#������8�.��B�8]�h�MR����*���0���.r�ܔCAqz�Z���z��g�,[wY|g�(�U_��* dܸ���>���mcy.%V��+����?s���)�Ғ����0}��G��yO���E��\3V��zҦVZ7��f���V��}2����
��������u��.�
���HX�
��F<�t��|���BIm$6�t�"�?��Ms�:������W�G�3r��14��(g�kH�+��Wk^�*l��?�{��3��X���n�ct�y�ON>�O��EO��R�;Ғna!Mǐɍs���c1
��{JI�G���k�K�I���"�����~?Q�5���J�����e��'.ߤ��i�O��� �?92� ]����}���_�Sx]��0�#Ht����П��`���϶�^�5��[xL<i�yj)cu�p�L���݈j0]���j;$�����w�?(��|�]aSl�ȣ�Ba7���ԧ'���3��`'���V�j�Y��c�*y"��qw3��+�������ޮBA��ŅBt_i9hF3g�תʄ�	%_I�?�����<,���[ە�0ბ %�E^l&�}�ph�J���2�YG������^�<ˣeL&R�_k�o���c9��vC���f��x���LBZ;���D<7�J�ߏT[�6�Gm���8T��T�����R(�h��G�7><,����䄻�ў�mg?�@%n�4�zL�Ov���D.v%�~�4og�w��6�.2G�p�B��uS����1�T;��������ӜY�ڸ��5�X��Q
��^�d�)���x7n�K����(�Бi̬�/����L�m��yBɍt� ��&�� �;���d�%�VӚDq���O�Ϣ�}�ISk��K�JH>�]B��U-��!��٭�&>�1O�Q���.�����CC	��C�	X��D�f�EG��� B��87z�V��W�D��x��9p�a��rӇ�2�9N����6�����Oψ����|`r?�x���+C
T�S3}d�{�����3�8ZZ&?s�q��"��u���{���g9OTym񘛸����2�I@65,��^��[R�]n���Z�'��;��u���b��qد�����8� �
�aL��L��g��̱�o����{�����[�<U�"�B���/l����	}��_Iy\�?�{�;_�����--A�Z�u����yb�m��0M\ ��p�^���	�4�vDv�{Sڲ�n�xLs�8`�qS�UR����T��Q��̟�U,h�7�Θ�̹[O?�Z�Z��3(�"fwoDm�����xǡ�m�h����X�a�8OS�	?�����K'���;�|t{�gp�e���c�uXW���)��l�z��p����I�}\�1�=k�uʤ�04���m��%�
�*u��1q+UE�s�'p�^Wn=�������`/��fEl���xuE_��,E��w�`�4n�2_�4g�>���P�ڥDg��i��R]�*nT����o"+�u�f����H��@��ل�Z���F��v5�v�H���1sB�Q�1��V}s��Қ�׵㭹z5^����\�#k��e���ȩ@��}8�f�I�"fF���������+�[�n_�;},�`�����KEj�O 4z�*<���X�A���झ�ݝ{��ÂO ��F�KaOY>3���>��5����QBb���AQj^����ޣn����l�z����L`N;��U�KĢ�k�
���Ku��RT�g�)͏�!��i޾�sT�O'��#��G#����i
O��7�@5�N[�)�v���=���On5{n&N��R�}Pי��=&A�7�ϭ���#�H�|�f�N�I&@�T�����
7��D���fĴ�_)G���w���������jrk����9r�RP�IWQ�HD�(�!���L�  ]�=jh�A�H-!t1�B�y8缳������o֚�<���.�u������PQ�
7g��D�������B�_g��j[��qB���!�5y�/�g�U�P�˃��[4�����Y����ṯ��F�X3D�����n��e*V��l���!�<<'C}�fg%� ����� p� �P��^�B)j�?��\��\������|����n�{чK�Ȑ����x�Jն*$������rG��̢z�8�Qmk�{�9vj�sY��k�Վ}����o��U�Ϲ`1/��<�Fv�W�cY���ܹ�������>~���e<W�~�`�^=�U=�W�D�M�;3���*� �x��K_��C�4������uӧ(�6o�zf29�6֎膿�� �9��M�z`�!#�9�������}B՚��,C���Q���c��)|c���}ҫ�g��U�Q�9^C]/R�U�������s�ŎUx��r���pG�A�������w��ß�~g��vLTF�y���5²!��-6�b���1���x�&p\�I�{�^�_x�?��t돤�҅H��H��~�wl�|vU>�9�k���xB����e�'4<���7vҵ|3ɸs_���w|��W�#�UM�l��Jl��Q�	��wi��x�u?�L<Z���6�'���"�Lx�D��Q�`KˇO�!,�X�>h}_��LC�j�ّ�֑Y�$(��!���t�"*��_��SPyֹ3���f�.���;əp@LWfݪ��0p7�u��撥�Wf�Y�aN��X�]܀V�F�4,9�?�
�.�d{����&����i���Q�M�U܄M ���Ym>�W?����9�Ӵ�k]��u�7�J�0��"'~$X��t��K�V}�JR���]b�2�3��Jd:g���r���k�d]��Ĕ�ڎ�wͽ�k��n@��b_���w �W��×1 p������M�������GL� ����t@-���{j|!���e�\�8�48�����Քj�<�/,Y�K��r�̖tz$�H4���L�����M�+`"�����S;�4����ؤ���4٩8�k�&����ڈ`����@6���3����s��[WDl�ȝ3l���t�8�o&��Lt��Pa羥Z˕A�H��N:u���\ bS����v�͎�>����ۏr�U2��R%o���d�b��czS�U�ě1�L����b�r*u���c� ��%�q�!
�٬AGB4YU�t�4�RZMw�j	ݻ�"G?��2|�����Z��XblǺܝ|���I�-�9������8��ae���m�^D�=�q�a9{�/'x$6t��5��Лte5\���o�!g�[ف����Gt�ֵ¯0�g�h�o���ܙ1�;[���{!9a��y7��+E�/�eG��, [U�V6y&�J�Mc�eOՐ}̋��Y!2GBE��^&�]u�m�a�7 �/��]�5��8���m�4�� ���������e￤���a���c)�Y	
�O��du��S �΍KI�uA)�y�P���^��S�VqZ���l[�&�:�j��T�,�$���5IH���9p���g��me�r�]aW�y���Qq�͝R�U/��T��|_���q��\?�'y�VZTl�,)*q���.�����yK0F�����`4�I�@~�s<�
���2Z���Um���0!ſ8����!Yo_��"��`OQ��D��g��h��.�4R.1~�t�ė1V��nݕP}�9z��)xI'�"GĨ��"h5��Ǩ@�[�z��$�d5`�Ĝ~��ͫX����ʇ١�������S�A��6��&��}�}z��A8ܣ�D1˛����q� �M�S�ZFV��ؾ��%�b%��6:+7��`�o��Z �	�.�y�U!~��D�ݵz_�������7�8�Q�����]m�ryq�e���gu+�	 (d\�F��u������K�����ɵD�m�S�6y$���I�Y����P�6`��}ӷ�k=�c����]�/|���Td*�"8�}�I���*/��,[�"l�槅3����o�",c��#m(��l0��(ON��C5���ww-�}�{�ez{(��wX.1���	\��LXU""�#�oʇ��x���b����W> �/wa+r�K�4b�ןD�m��:J���MP�m������7�Gه��N��T��#e=C���Z)��&_4jX/�Y��3�l�z��r����V��E?�~&���y-R
������)�q�
�0*`j~��/�q��LZ����&4Mp&��gi�n��!M���/�"�l�[̺2�ݷc�)?��P+�q����h�S������j&�o��{l��ec:,��ߔX�����AK�6���rG[�?Lq^P@��m�Ȅ��ލlEo�fb޸�)hi��ƪ�7�ݚ��gn�Z) yHk�_������X�E��_���s{ a_%�T`׳W5?Z}.�C;xD�x����^��ʀ���8�!�CV=~j��EJ�]Aw;����~�]�F�����>�vq�1� HEHY%V5�z�P혡�Y�|�^}?PӍ5ISpU���ѵ�6E_j]��͚���-
�Pu�u=1�3�m@Ц�WWn-Mx|��"�7_��y��ј�DU6���N�Ho�m�����q�>�Y�c�6�ޒ�t���w��4�1�K��f��zӸ���@˴�۩2�?��@im�Sj����Yr��c�D��T�by8�(��?��q�:�!�˾��42��TSҔ8�cI{�P0k����_� �M�H�
�g7l%Q��jw��:Y[�.<%�j��"kSd,%�6D\F��S��h���e5�}k	���3�i����S��HA����fϰ9àt�y㣭��"�89���:kn_;)k�s�<�紷O�(nbV!�̖�*�E�"� *����i�6O���o��D��4H<�.N�޹��ؠ.��e�N˵�F1J�1O.�_�U& 2)Fc��(�бґ�1 ��3��fF���$���d�������gJl �t�h�/ݴ�O�,sPvz�'/{�������U�ݠ�H��A8��P���8���)K�{��i8i��Ȃ��6s�AZ�u�#X�7����J-Q�Ɨ{U~���v'!z�n ����I���*B�i� y _�&)�G��/U��cs}�S�∴o4�5	,�R�\!}Z ��^��u�����h�I��X������h��4��H���gW�on'9�GHH�+gv�"S��J�{��l?�YM]�]	��&ܱ����������#�:�r���:�e��R�P*�zU���5��OV�g���jZ] ��F[�rFv�7�,���-��KM����%��5 �
���K~_��ji��F��F�q�jW~�c��G#r�q�g��%�e��A������`�i�
�s�]�`X�t~������ss� �q')�*�j�~z�,%%S%��^5���.5�+�`}+����V�~�G��vXJ����L�$2<)��k�>�t�2�����ͥ\i�#4|z�^<R�8*�n��l��]�U�1,�l���Q�̠{Òr�Gkבw���u�
a��b����R4��̪�.��8�*�h�7���L����q@���G>��ןt�a�W���9�'�oC�E{F	Hx2��:���_���RH�rW�j����Z���O>V�\
�q��_�=�.x��*{=?��0����[W��5�9���H:N�BR�1�ɪ�j�cb�+�y A��t�9���U
 0Y?Z��h���m� o_���� қkv�����GK��1�ha�3Ո�jK�������u]�e��s���y�t��Lx��(���ˏ�,D�rܪ,O'?>�si �3UE5�&���~G8��a5��4�ޠG�Gq�:���˶V՜��Դ�G�����'S����X�����2`T��^6��~���=qK;}���Yg�u���3T-UM+��9h��|e����n���A���|-��m�;�Í�����9��l�M�����x��ԟF�h�r�M��/�p!�19?�^)*��b?�(.
8{����U���<5|+��x���덵�I�VX��@����dSz�����ኀx���A�j1�z. (`�>X~_E>e5cI$֋b]�b9MՑD��n9l>��� �t��AQ���r�W��	��o��.%�k���]�m��ț��Q$��������<����w�e]|K�Ҋ&e�՟�^}}���5�,F�rUHVm6>g�8�ԑ �t_�U�[�H��5|��6F�5�I�p@�y�/�ʗ0��G����8G��n6/U�FW���S�&(	��1 �YTX��L�ϝ7� ����1n�Yt�A����#f�p.q���;!��AiOȀ��ٷ>�,�5�s�5WxT�Z+?�=�B2�R��:�؝)u��o�}�)�;��z�-�/caN�]��� ��(a��]�Q7��5�%�2�8|��Qz���<�SvV%�:Xp/wk^�4�XwE[��!5�O�>}23��,�.�;����/��!���\o��hm`�Q��)����uN�u,�d�GެdH���|T񷃇7�`A.�������4)@�}�ʣ���G	�K	a�ϼ��r�9�8-*
����{Du9~2�{����L8��}�H
>?��t�ݣ?���������C�$1;��t�cS��@��puiO��B,�f���D��YP�-�aIY��xJ�5)^.S6�Z�8�S��;��^;��t"�<�M]��"Fȗ@��A+mΨ�_��9��5z+}�����˾�c/��:�w��D�e��r��-�䉷���{8@�}�ٓ�fT�LͭbZA9���	s-�Vl@���I3:Py�����w���Uu�HGX:��ݤD�T���j�@��k�Ҧ�ܠ����Z���C�9�vD�Ļ�S�=8W|����<��J�p������gN������~���M�^4
Z��j�4J4Xo�����f�7F��߭�;�8������	p��&ݪ�Uό��Z ?-��[�i2�=0�d����#:@:L`������&iӤ�O"�nk�$��+�gm;����0(\�I	[{;����2L�9�b0b��<3wm�Xm��	���8��� `��1���8���z���F��i�MjYH5�G��j=��J�7",����-,�ļ�ӌji�%�,!n��XTc����F��ru� zg�*Lb�#Ζ:+��!g�W3%bVu{�T/�d�/:�S���Y�E@��
�.4�����mJ�iI�Y� f��
^��+�6ؖх֛�b��]Z���$�(��n���(���ͫ^nZ���\�G���=��ńU|�l�{�`յ�}�"��̞�gV�8�{�k/�8��6�02���y-�$�'�a�V|.#5��֥�[u�q�%�FP��d�^�y��q�;�Q�0��?&��D_
8��'~��Z#qc!f`|U��&rasƀ��BC��K�'�ۚ��f��N�Y���4�Go��7��Ü�k�o����p@w	���6��ix�nwF�i�ـ�Z ��Htf�>�I����ގʻb%�����
��9�%�#����ez��I�u򨆋]��}  iK��6q�y�4R�Y[���հ�<�����1l`���8�-��!v���I�����CG�v�҈\]���|-��f��am����o�B��
��]��,˻w�W��՚���M�r7(4����-	Q�_>ӡֹ����GNq��;�T�����w�����T�;1�!��Fak���4��L4��U��m�H:���.b?���-��fK�3<{sĮ)�>p���^��'.j��xwb���
��k�á\�i��[�
�|
u��qaW�H�B��q�t�m��Etx�pdk��ڼ�X�h^�u��	��#�x����QK|��J]t}Q�l��a���=�^w�_����J����C*;� ��[�3>d�k���p:�c�W�E�Q��ǋ^z9&���T�nHF�u$�(�)xk����ҫ��������UO��pY�.�����o0��%C��{+�p��n�TV���7��l�Í!?1�$�׎�ey>T�S&�7Y�>�%o_&_d�K=�z��S��Q�y>$f���kw�9��}41�A"G#�1����:�4J��z��烏��������gyM��� ���8'�l�r���e��<�N�>?FI��2��
��/|3<3����TZ���p�Ƞ��B�2"�Mػ�X�3�љ��Y�h�?'ez�kpa��� �bgA+Ymj=�6��^=�O ����.�k�??z��F�-���0SY[�jg�}��ѥ�gU�����&�P�+�~�Z�Dv@��=���K}Pc�B�����Ŗ��{mˤ���O�7h�	���f7�3 |���V�(�O��%���˛N���=�����~!�B>�)�,����4�!-d-�rc3�Aߥ���)��r���_Ы��Xg�}p�˷W�EFE!�_�����<`��^#PVu8�<��T������i��3�4�9���Zqŋ���L�9�vHi�!Þ���Ĳ	�<^jC�4
�9S���Ɇ`�����7���@�߿�����j׌�CCr��w��B�q���+�}�Ϻ2��<	,��)[�⡲Gk����k��s�XD��J��X�\���P��"�w��k��pD�/�uE����?TR�ȇ�߷�{~��p�	8`N��� �o�b�ƍ����u���]�jG�z��v@P�][�~���`�B����%v�`��+�x����t^5�k{c�ng�e��k�$��4V[���K��I.o�<�	���(J���.�/�IA�b�΍��e��,޲��t��Q["��\��?�b�'�{��4JD:���&}�vr/�V$��l�i��4/����OZ���}q�k�l��[2�	-�%$�1�w�6`���uo��
��g�q�- ��ȁu�KM�үF�k7���3Gk���O�MT�h�p+��?���?Q�D-ts9�5�'v$�s�;�dἥ��>uc��߄�G�H����O��q��Y��.v$z17�'���E�/Yug!���
f�`i?���bop��[��9"Uoc�GWp���}��ڢ6,�Pw���ٵ3�(�.~#���݈/�o��V�����2l=ve��I���x�4+���9�M�?}�ґMoZj��|�Y���+�� -�Z��n@ ?���q�^oC�b9VUzf��\������������B =t����b�S~Z�yqFƓy�������ϑu���O�:�O�Q&Q�<~}�?4ĩwڄ�zo�/_��O��|ރGm���͑�ʏ�C,�����ٛ��܉�^��ޠ��g/]zP� � �㠂���_�;Q퉒R�ݮ���R�	{��Kμ9�q[�Yx[�/�W�����Aq���+�o��4��;5}��222	�����յIxg������6K��GQ��q�3M=ٓkfY��^m��\�x��F�\���䵽y%��J����,Ǳ�����,Q6ɵ>��E��<���E1���|&�p"���|22WE�8�8�ۤ޲^y�x��K�|�m�t��Ƃ:3CR�<����������"���JC�P��pxc��aj�<{d�*���#��0*�s(8��u��y:M� I���mK��=o*�Z ���0��v����&1�m��6
��K�4�������
D�y�T2���n6?��Og���;h���\�����%�0�leصk�g�|ʎC q38,W�<�y��]�~���:'{�pE& J�� wB$=��(�������)vw�g�̌U ��^�2�+q8q� j��G�o��c���W]ʱ��gv!M��;��W�(�x��Z�L94����y�Ov�E9���'�׋���w݇��J�����B����A�-X� ��iɑJ�֝X���c�nk1;�-]����㋡	n��B���E_/�!��Ԟn�Ihf�M.	 � �>(�ݕHP<Lq��͐���7|c�s���"�����U�o]�^���$� ���3=n5�L�`��#��+�oTX���E�%)��P4NV�%{[.�o�=��'�6�oE��R#vC��C"�\���0JS�8�K���
�O��f�y`Hy�����^��&n�g�_癮��IՋ��y�(.z��\6*���Lz	��=��m�2<@&�9? ���51�i�ݔ�k�6�1��Z '�脮�M���.�<��i���47�a[���5�<�C�9حI�ەh�3�� �� +9C ��۫=Q�0{?���&��3I�V��[��#8��g�@6��*6�Z�'2Zqۋ��	11`�}��i/?m�^���Gv�̍���{����0f�U��-���f*:�(�Hr,ȇ��ùb�,��L�P9p��Rpu�/"���L\�έ۷ۜ;'_�@o�@��{��fl$/"E�t��~�^7��*`#�J
_���Ͼ��P�G�e�l.D/�~I��މ���<Wp��M���I��eO2,�ee":��ζ�v"$w��J8c��!K��Ke�!��?	�g���E�Ԭ�@�>��w�R�su��)�פ��\��&%K���~�[��+KA���l o:���k^ `�,:�(�JP��`��{�X�t�w�9�7G:��(AZ��l���[kY>Һ�Uqq�1%D�����_�����i���
�.C���׼���Y�&W��B�:|� A�X�4m�:us:=pqC�8+G�^��t�y�s�7F5������m@9o���۹g�z~�kgkx�Yu�ʽ�ۍ7Ϭ�I){�Q\5��r�ح�}���4SM�^���;�e����E���fi���f8�z?�	��=Z�D<z���YJ�s�����໒,@��7/��UD���+ N�{V�]��r����/}Ț�Id#��?o�ޓ�s]��O�u��V��:���@�*��S��	�,=��f�G"����p�p���˃�X���"����=EM��~�/C��~8J�����Fk�u3�#��x�3Tl�DP�w���"ӅW��s��pĭ�ij�^5��%b?�/��1v��C	)0�ƒ3|[ůP���#�&��.aC;���;��s�k�3��m[#PƐ�Ə��UٯV�>�ǘ?�d���/̣�2�u���1��[^'�>����`|��^��-���v5Z�k>�3��>�����'&�2�b5g���3��c�)m�Dq� ��W�ϫ�kl|���6��-С^֍��[w
kIA��|�`1R't�#8z���H>�#��o�Z3vL�����7�BXz5�1���ꍲ|��hH��o��i
P/��wN��������3cf�����T�o���
�?۬�5?�t�)V�1*d->��
�g����z?:�59!��N�>�{�k�۟o�`�O*�|:�
@>���K���_�������/RJ(���h����@.����ɡ��6V���G[���(P�����t ���^����h�|�������e�/�5��Ĝ��*{]����/�돏,p��c�N����BZ�S�k����'vDT�Xy~�I*��v�晀@;�H�MR�t}U��'&"-L#�����(!} ,vy�q���Q� �q��h��g�X�N�ȉ�j�C_��n����Z���*e�G����g_���O�\Їz��>P
�R�Kw���|D��ˣ�j&@L���V��;�4� �� �+^|�J��+��$9KGwA�F[�����H�y��m]�1M:v�p4��zg���̗6���@�㒳{ ��*^�H�,;hr����7톮�?9��!`�nI��<��sl0B�CL��̴�2�xDO��'(H��=�A�۫�dZCD�]�ؕ0��3!����N ��
��9�d^���`�� !ngJ�㈊��<� ��ѝ�A����t��F=�k�I;Ӣ*�&��ՅL�D�ѫTi�<[vo�I�w�lk\<����}4�b%� B�ϢA>�}>]>��ي໨਌z`d�f)"0����͹g-���I�:_�9=
��}���^kF%}��~�E}����CXp�п'5�@��\�(<k�n�D(h��<F����a���E�
	���|N趨%�8���& :{�A��G�o��FN���BYYd�^,>ܑL�j�w-� �VV�uacy��|/Lb���3!�95��4Z���>�������,o �kK�8���$�vS��a�9<U�����ĉ#&�����*�o���TE�QU���(��{�pGV�돇bm�*,%wg�ʛϚ�������M�]�"��O3�{�TUZ�����i��n_"�֭�a��$px8�O��]-�.���3��C���\�N	�����w�}(��^������x���&=��5Bp4<��ic�!a�#�]S�Z*4t�L�Ƭ+���kJ�xf��­�@��Y7�o�����iQHb�~�%t�M&�Ĉt&�܁�LD�}��>Nm�p���ަ�����Z@�I\���׬r��ol�>�l5|�_�D����^�|>���Ϥ��P�K6:<�>XTF�ȶ��蠖i��W�M��r%l�����]� |�wV�߈����Wb?��35�&���.�7�7n�~�S���de���
��_��If��i?z�p�R��~1h}?��T�`���TO.ع=������W<Zh?d�7��s�)�����k+������dfߛDf���d�h�8��
�zZ����u7i1���/�F��c��v;�Ҟ�b�/k� g���[��xK���b��L$���MwX�1�#>��ZZ*��cb	%�'v�)l/ ������B�\�� 4���i�0KÖ�K���V=9*>��ox��6C�.�$-F��E�h>�M֚�%����	��#=ާ�F����P����{&��-:RcDSρ䕼Z�K���XK�`.�n{TU�w���p��^Auo�eCC��5�,b-�q�?GGN�̴��:�n�~���� /�Z���p7����'��8R����(Bt�=��m:��-��8G�(c~��ΧP��+3Ϻ�'�1.���ބ�'��=d4���!��sTܶ�q@���NsJ�/ο��g^.������(� �49pQ�>l@Eb�n�;�O�GT�bw�n��2VѸ�ʤ�K݅��큄=�{�p�����.aъV���d�`�4��0 �j������N�Z��~�pʃ;иZ�nv>����_��' � s�:����� ��y99m�=n�1'�"5S�ܓ��k,��k�h�������}t=Gg5����\�ݔH�}��ڥ���C�Ҕ��*�5w[J�~��n�����v�^����S=�0�'�����dA�Yh���^�i�� ��M�2�M�隋�y��g����U��l+��V�$v�^���*b��5�~�Z�7̻��a��~�ޅ�|X�i�j�>3�����Ȓ�冧{r��ε�&��#$�`�A��s𨜐�!H�T:�uRv�RnU�LPS�]�"�=�PqH�Q�,�Š�7p�M�:�W*\���P #o���Ѱsd�o�!����N^��h������Oȇy�/4���Qe�qp�(��Vo:�d���oH���&[�����U������W���c�LU��Fm�혟8=��(��;o�5�	j2�ʩ�{1��~{)�l6g~E*���C�������K�9u����f�&��mmU׀��{F3�n�"M�$vVZ��! ����=�|+�n�O��Ζ*-�U`���`����j%�$]O�{��r�R�$m�EORC����|$p�Jw�����ɞ*������ZC��D���m�Js�֗��Nm�j�>����äT�	H���Bp$S|��+�VZ�Qx�BI4�ɶ�AHX���*�^�7Q%O�Ы��͙<y6���*����i�յ:f��^<����z��0a���P�īU@;��O]���ҍ����������M;_��-���s �؝�>�'��U�=a�S!)��Dr�`Ee��c��qg��!�ى�x#}��E�#�Q�g��:��&�w�>/�}���W r�U�����s���>F����w��O�m[��]%|����k�A5>R$7dmm5��o��� �`d�ut:1p�JNM'��c;x4��1n�6s����vG�ٯ��9�d4Pw����಍�9���uO=��+�.���?�?�&��z��&�Sw������">qh�}RRd]�IsJ�e�*�PQ�k����e����Q��ܑ�ͫ��嶽u��/N4�Y�f>I����]�'��3FsF�4([M�އY΋�����ʂz�rrڑKkkT�:%Q�;^ȫ�d����؆��ѣ�a�U�l�O�8:��𶢚��S���r�5�Н`K�p�Z\�NE�=��PG��w�D�2�I�nfb���vp����p43���Zެ����&���oM�Y�v?^����d`��h�g���/���(U�nU#�:�O�[�+8al�&�����׫�M8�������ƞ��/T�m�� b�]���'��o;Ѷ�	���-Z��D���S+e#_><�t���u¢J�6#/p�zV(8Y7+~�oS4��}��]Vu�3�d̵)�VTTx���v�������j:��Od�V�;ۛ��!��n Q��.f�uߓ���}��}��Ķm��5Bz:��̲��L����rh�!�:����"R�O9E8\��t$2�~ Ҹ2��Ϳn	���ZG��7�����b�:rX�G��PJ��!	��;ã�oQ��g�z��]�* �?�&��%L}+y����[�w�D�u(�Rϭ��z;�L/�o|6�`xhb1g�\�|5l��|��}��ݶ6䤼(� $������^����v?M�3��Dv�+��g�����g#��%W<�� PK   F�X+���  D�  /   images/5cebb09a-e86f-4cb2-800e-22da09d26481.png�yTSW7k+u Z�	�5�����dK+�т*�"�2$�!L�
���QF��bŀ"�@ ��IH��D÷Ͻqx�����w��ֳl�9g����>7湴��Dz��EA���k�6�������o��*���>?���=�'|^H�{؇@��A��W{j�<\s�W۳6d׳�c�.*��v������E���/�_K l �~�i�����n?=~�d��y�>����g{�.߱�k?����n��������k=.����yAʶ�S?7/ot�Qi�y�u�̿�]1�����_y�͜�~��z;f��ln��	�	��To��*���w�y{YJ��|���\�wr�k�0�g��2)��@�0��P7`2E��]��Su����\�64��b�BU�c�C�qs7E
{�U����|�
d� d��\�դ<M>��ᖼ# ,��m���/;K�5������k*�pnyv����ßM�GV�m�o����߆�6����m��m�����	�(e֚�ܩ�wW�^d�����RX6�,H$}� �o�h��x���X��p͎�Q���cNKCnBI�q�=qHi�e�{O�1=
x�k��U���m�n�$[G��3(��S����(WX�}�O��	��@p�9r_�6���9m|!�X!?��5>B?k��9���<W{���z��˿`��o�_� �ix�2������{�7��k��{����W��r����BE�z���V���7/��e:�I�ېc��2�?�)N�oL	G

�������/�O����"���<�Ot�"�<��,�z瓂]ǿ�ϡ.K��l�V)�8K>/��i|bH�	��w���*���w\ &�[��F��Ld��4�2��f@O���Ӛ�h^�d�+��K�������	(��S�|M��;) ������F�gAB2/	?��{��8y��v�BX�-���"]CY�����i{�\���D�=��j0���f�/q��!������M�u��>��)I�d��dK�nɁ_����Xދ�9s-0`�R�c8�@@�5����5�/$P�]�ر� �tZ�J�+R*9��|@\��5��v?��>���:��:���$2����Lb�z\G9��~\��.'�ny��!��-�q1Ș|B���_]$���	������|oS X&p�mW�c��~�?���{@�9�(���uX�MH�-�0P
����`����$/�������1��1F ����7r)D�v�s��Z|;�\h�D,1W8���gƚ���8f|��J���W���~!Řn�ŵu<��K|���ޔN�]�.�v-��r��7mrue�'q��L)R��+��¥�����z��ϑ�g҄DM�f*�r�Trܒ"S�+�#�+����ϝ��f!(7@?���9�#�?�}�+�a��כ�+��EL��\��&�I��}����I��]��g\B��Xe������)=PI�Bc��<�p��Kb�DB|~_��[$� �Q��=��g�����I2�uC����,�=0�����霫�3h�����tG��n��!�Y�^�&��~��"}d�}vxf�=<���:�G� 1��3���`�}n�ϴu+/?_��nF�޵��D��x9��k��K�n�i��+�0qa��1�y�8��h5Wb�م$59��C4����.��9��ӀT'ɛ�<�T�/�'6����~�򼚄��)�YT�\�	���)���/(�Ye�� ~��J]��*����-M��3H1�nlش-�{	0�`{7i�$�d陼'��K��R����ԣ�����]�QG��P.N���2��;��/��~%�mRN?f��
���<�WE�s-t 
��v�Q�`��m���4@FfUyrv?�m�))������-�����2.nxJ�Ǟ��߀^OJ���X4F�M 
�m%	maz��k�j���O��� l��fI_6.;�G)E=ΫM���/N���쳰,F�Z �z؅�n��?؁��< ��S���¤�h��Ge l4������,�nY)����i���8���>c�7����x&|Ό~LNߖU\��*��9.�S��(�5����^����@�Wǯ�*�Pq��R��ySL
����oâ�z�T@�� �ǯk�.�)�kD�G�e4o�����o���UT%+?5�DO�/�pƁ4����}��"�sS�b,�B5�/X�ٛ@Gr��!y�6��ē�M8�7�I U��� ��[Z��B+j��t�|�2s��R��I����;v���Eʢ:d��ЙT��ob���l�}/!�0�_P�u�[��gߊ2Fu�܂Y��.�T�����f�>�g�?�nY�������g��Q���D��R}=ax(�^~��?06����G/�v����p}�37���o�����s�"e��X�����z�l��cZ/�)<�u,D�Sܮ�E$ �CWL��U{��� DC/@���PcA3��$Z��{7�(����a�]*'��� ��̛FP	�g�G��S]D#=�
}V��.=�칵oL�\gɤ��Ìl2ܚ��N���i��6@KI��7U�>W��ʷ=�i]����Y�ݓM��[�{���ީ˕�ח�>H�=/@��kg��4�|*πTYU/n2
9��֕��^H����.̥OL��&�I���{����]��Ш��k�y[���X���d*���D؆-.*��}�l�U� ���Q����l�e��e,?��b]D~^60V��4���Ӏa�̟�SB���py1�OT�78���-ߎ�5����Dx~ء�,>@�jeSҼ���������rt*�s�!�[ͧΊ/S�F��x2�A�G9P�GT�� ˞��@���'��F�L�W1�u�p�X��YAR[,��8'�$ 2����0��o�=�
		Z�/�dvWC�O���{���.Y�4w<Yw� �Ke[�v����˝���Y�Lw��^��5oW[����e� 5����a���r�/��Rq/��.!�kV�����#��W7�h����S��k�|�Ю���)V����<+KbP��i�,2t�=7�����,g�r�S�4�՝j؝�&���X{L��^�͝�H�����浺K��,=t����O=��`=�k�i3A��xM�t�y��W��^�����O�gﱦ&��~M�pG�3a��f@3H��qo�[΁���ﾡOm%�Z���53�9o�,E�aXĿ/����Bx�_f��;>�B6����M-'�x(���];��k6*3�y��"�ץպ^��r��r8e:��M��%��G�F��E�Yӯ&گ����/�Uk�_祻����}I��hi���2o��6�^��_7U0���p�<��%�?LD����л����g(������ ~O�./o?r�}��y�3��Z:V	B6��U��3A�u��ʨd�jD���\�Κ����ӓGv��n$�[�l�} Ȉ��H�H�m�O[ó�3MI�n�Y~X�������F�A�	5�h*���U�k*�B+�7�Ŕ�(����YY�ɩL8d*Æ9ߦ}Z0A�O���N�'���r���Y9S��wnC+q�������2�>��N��R�5y{!wK��(��x�Ӏut6�^�d�_&őo;S�M�wQ���}傘ۗ�v��?�����=�2�ϛ�J2A<�#��nV�x�[��� ���]�9�]��z���,�:���Llʖ;��� T��3&�_����^T����2ET��q��N����9}�O$�[��v� �͕�,Q�̶?��܂�Qp.��8��uE�B�%5�X��nb�W��j���MY�"���U?~ j'�rA����p��&�7��,�0�Χ�K�P��sE~�*�ơ��r����ͬ�?�Q�i7��̏��:8�H�2�9/l�(H<����^��#�$;�G�z\���,��t��իޗTV5���^���l���|ϝ1����v3�[�9+�je�ŕAc��hk��R�����'@�h���FM��m�	[�b��`��baW�a=�((��2�or'�T�9�pZ����]X��,+.ˍs@+�{e
V�K�n�J�5(�0��P�$K�Գ4z�����wK��nO,!,�N����k��SE�j_��ƞ����z20�kT�l�3������}�{���R�A/=&n�b}�k���8����f��YŎ��DU�?��n�����䐻~ؘR� �j�[e4�;:�ye$"�C�w(R�3�o��9���{���=��:�6"��x��
k3������Ṗ�ɑ#p���ͫ���?12�^m���'t��2A�f1��Rf�M��h�	�D�:[�����h�:���p��>E�JuY�p�*Cʇ��;�`JLz�4�e:2������˗Fb<�f��+��J�W�UG%'����j�����Âq�l�_�τt��@ς4�A�5��|߄�v����61��Ϲ+7�[�,���Ώ.�����}5XA�)�X���ޖ��4TMWу��d�2?3.� j�!�9���~+n���rM�MG�#Z$/�¢	cd��6�}�d	��ȟSd:1��l3fN� �d*O�B�f�sC��g��<�}�=�����^��Ct���]�'��$d'�IcZ�3�ӧ鑓��nر��؊@*��i�5YyrJ.]�2$��1?��WJ6��C�xoz�qxO��-^�˭^>���U��d2�!��ݿ��5�i�իF�'��:�fBWE�撈����s#6s��:!�Xh���R�!4o����I�g��5���޾oW��"�����(>��F��=,O&��
�ݱ9��4(�t6���8��kO��}��l�뚖���B�T�@�I�|�>}d*�HUd9*�9�p�ԂE����7�^>�z�u��m7�7��;8��ksD��%����B�Cy�90�0ϲd<ռ�X��A�3�v>{��1�aEw$=�%&�S�o�:mW�b�:zs�LNc��j+����c��e��O@H�Xi�8��c� �W�$g�9�#����1÷o��&r�A�.��j��=g��MV�tSjy����ѼC�F�/�b�Q�W�@��Gy�"�Vrzώ��Y���*�6]#V�a�G���nP�^熯fl�(ǻ %��!`K�����"�{jd�Zw�8��xr�����
,����?�ԓho�F�rwc�4�c��Lb+��F�P0�[��2�P������M�����>z��|�N)OJ�eM����7�E!v�6�S�̕�#�;�/�q��쌺��}��Y�v,p�W�d�R��F��x�_�V8+Qm�WD��>X�*�wI��R��\ϭ�}𺎌c�Mu��2��c���n�L�;�������HQ�Ik�mS������ғ��*O������:���d�oE� �OǷ��'?�gd2��[�^���3�*i��lk�G���F�҃S�\�G�L��&�ۻ��u) v��h��f��+�T�����o�"F�_�ʤO�	AP�v����<�9:�wk���K�=�X���@�ުN��{��`X+JP5���ϳ���F�9?�U��a�4�R��m���f2P��Aek�0]�"z?�8��044����t��s���93�}��'bz��!NB��[e�zN���X��7"߂NaY�I*�Vj�c��i38������0�ct*���4��s�J��a�ݮsq��'��}�3���vO����C�BJH�LIP1�*OO��ARt�oc�յg&��X�EO��}����%C��dD�Xi�ዪI�|�lK�ڷg�sĺW�1���S,�xk ,X���,c�ޥŦ�c��K��=����a�}���4Y�v���T��2>��7�KX�iD�
NV��ED��02S#u=�*���Ao5���� :9�/t�����u������}K/��5��y���U�L�mt�>�K�5��'ℸ�N4'3uYc�d�г��H�rAv����9G�0�
y6�he���:��l�Z���?l�\��1�R�a'õ�(�������-WD8��̅�8p�s����dQ��-���G(����5o�����Qf��]n�"��p�7q��:g�H���?YK4i���]�4dQ�ץ��U1<��;�G@�d�x�_�6_M���'�V���r�e�����_���#_,�i���5�N��YGWR��?�O�ׁIVeW�9F�s�<mo�#\���&e��p�W�^���ź8�5��כ���CR+$���k��y��nWx�p��S�i�����7n���A�g�X�{���g��5j�����C��	")x���H$���[+%됐M����i]�%�q�j�>iꭠsނ�<��HV��OY�f�#$d,H�} On���Y��� ;g����U�ae�,�A�"�I��՝���"��ꉋD^�6�;�_zeF*��r� ���P�9�{��� L�F�$�h	�G�N/VH������%��I�^A� ь3>%9���^�;��&D(O^Ȓ�����x�,%iis�������?�elb�5Z`�]]u�[�k�N4�YwR�I�k6�Yp�C�%����$"i�u�����G��?��ҷ[lւW|���. ����Y)G�6�w�/��>�b��5�1�k��IY�#�svA3��~3��5�'�3@�_�e��!�G����iI/�d�O�
�w���j5�	�~�����'B��:�g�gB�;�u+��+Wʽ����T��%����ol�q{!~n�E=Jv���(��۽tٗk�:Bo�^�~o�*"�mL�W ���l������z�0_��ܻC�̛!z�sn��iV�C$3�Q��!f�+ -�ˁ[�d�Y���|�FS����7�����Ր�>��vv[(�l��A)ØL*�]�������&��xRnC�"]N8�N#F/�;���d�,x�B��M��Mi����M5w���(�p����ղnR�뒧U�+yD���::|,Zv.�h�ic6ȱ��v/�(��z]7�����F�F�}N�U����A=ą�Xaӝ�J6������=d\�����-��W���x�]�A.�-�1��p��Fr��-n�0Hb�Ͻ���e=��XԀ�|+&+ł{84�<�6�Q>�#`�m�3g��l���G!�Q�U?�e]o��{���@��a�+�e�p�)	�L��ҋb�1c���0�<�'���=�I��뾥����;����^��U�ǖ@��U��О�,'q���k��t�J� � 6���r�v��6 �O�&�+lm� �lTvqb.�s���|�<�����"+�Y'���>�W\�o@��0Cu�[�d1����<������q0b�����-��?��Ϗ�E���
�W_���ui��(܅��"��]�n��
��Ћ(&�/5U}� ���?��Z�?��̙.jP7J�}3�x�ţ�طKlA��m6�9ѼK��d+��6l:k/��hE67ѝ�����QY+��6ő�_��MK��_e�_��Q���j,����+i��<"@>���P��R�t?<wφ��L|UkV�	Q�Fу$^# w沼]���CJ]�Qy�U�U�	�Tͱ�>f�=���J_���~�e�m����Q(��Л��å*#d�)�e��8q�7��[lϕV����b\���%�s �"���/�:L���B�ܣǏߓ��:xj��>��_�?���Ri2�W�&�|�֖<\H)0FGy*#p;�xq��TE?fj��$"�����#
L��|�et��4�
E�zص�f���;k�ʦ��yy@�a�����"��X��y6���	�,:9������̼��h^|83C*���'
Qc�˝ԃ<�S��W�Tp�d89JL���#sޯ�C��Y�G�_���C�Å{'���!g���Wa>PӒ[!7�Τk[�s��	Ǆ31ѣ�%� r�4"֖�%P}3�4wo�@!OzSn�t�?jۦ"��!`�U;�Hٺ,�r3'���y��6���k*�Ȑ����� �N�����o��*?��V�K����&���"2�>=2������x�ꂝ�:�'����T:Q���{�i�s���;!*�ź���2;;a�E�>8���tV(y���S�#�v�N-�Z�:�7O� ���E��I,�ԆUN>5��n�U�١��F�w�����s��Q�����'|�r��l 9\�=�]y�5�c=�YsK$�N��0��݋���ħkn���B"y�77W��ߘF��2
�,i�5ֆ�*���Z�*�<߄��0}�Rcc<=S��M_�c�y��U$�e��v�}�����4,�ϻ�ɒ�pB��c�u��+ƶcw�̀]oKQ��ȱOUQ��d�Б�/�5O�N��O�.V��ѯ���簯28�Ra�Lb��ֽ���W�d�*#2��+{�+h��u��g�!y#��;����h�#�Q̖4<׌
F.z-we�>�]D�)j[,2a�0S,�����"�8��������)t�;����8�	�J�ؤ'�{���84��{��4�X�:u}����@�7�`U�2[�7F/��/��,|�M缀�F"uK���x�Q���� @0�Ǭ���2K9��Tj*���V�{R�!�X���Y��{Fr�}������҂9��z����*m��'V�u&O���07C��`n3|Q�JOQI��L%�᧥t�~�H*`��Ah��~'�߃`0���Eu�Ƨ1��v��B�y�l� ���v������Ij��&���:��V �AV�D�P�Kb�2��z�"9$�����#�l����T����EZt��n�:�O�0h�W���\}!�W��*�mXA��@r�0������߻���,B߳��G��P��\�U��_���ܝQ�p���Q(�LuF�1];��'��WEK��M�u��� �o�Zՠ`��=tt�&-�o��w�k�b>��ԜPQ"�V��N����gY{��֧ؔ
ȧ�ﭜ��%�y�5�LNe޻Lbx�M����V��qs�������Ѯ�۫,�Xюcok�$/�����'s��3T�R��Nx��Z��<2w��һe4��G�᨜����JWE�z&o���ס������<u�-g~�S�w�D	�����'	(�Mb�2np8�x�v��@|fO��NM8�'�9�Ei����u�f�\u.���u����M�c0L��3���\�\��aw*��~&5�`��`&�X}Q�@��)�ܰ=�J�m�b/�-?�f$Ɇ�є�SYVg��5�V�Ƨ����	�����T��W���ط��9�^K��\����7q�L��TqWS�0�9��]��6��~f���/���t�"":��.I"�dl�[�J$��pd����q�b;��[O���&Z<׭���&���\�L<�\�>@ՓG��O�mﮬ,��7���Ń�r��L�mFb�X��n�+�L}:�e5��7]�]k��u��;��������78��M��A��(�~0������M\��׎WaZ��?�k�C����%�S�������j�\� �e.�A�ͷ�KN�^_�?�0�l,ۊ���?4l��;��s�������c�!ǖ>������W���46�d%%���6F�M�?�=�&��GJ��{�%���m� oY�+u��%�2���ލB���O��1/�,B~�8>V�ܡ�kVZ����y�I�jnk����!�Wu���Ti�l��nz��Z��UUAe|���T�iw1�����ޞ�&��G���@�W0OltUb^Pc�0�;̺���:#kC���ix�f@��&�um��1H��������$� `�&'CrP����	����4QPn��14;�1�<��w�;'�e�=�`��y-�����-�o7#� �\�r�i��b�� I��b����eD�W5��;9�s�����EF�GM�� ����#� �苩F���w�\%�����.�5	y-����l��i�B�(�YQ�� ;�c�����l�bu�ȿݾ��Ǯ���t׼W�s[o�m�J
���G�6��Z*���EZ�BάS�%%	N("�}gN���iCEW����J�O�c6��iK ��E-�����|�P?�H�%�$_ѺoH�w!w_�R5�!s�'��M�:�&��`�D���VG8�$��{ �'����B���W�.m��x��&�T�3�I��)�ÊHg�;>X��/�M�
��7���Wj�[����AE���`}�${���DG �����]��j,E"�����}:�R��ԡM8��w;X#������]�g�Jb%�:dٺ	E��� �V�e-������M����z�����WM"zl0�$����V(�~��!S-f"e]�q��Asl �}R'łO08ZJ1ʣ
���^�h�����!�*���#�s�-��R�o�껡O��1��BS`��i�Z7\W�,�h�(z;Y�/(B�V����D����~��O��^�C����Jt��H��`��^�UZ�����A�vrHE��:��*�Zl��=F��] ��r97
�{(��80�U����׬���2+UQ�,(�dGlpn��Q�^k��V����7�)���B��Ƭ}��0�I��L_qBṄӃ0�!]���Q��<��)c4J�\D�ښY��
�]��{��&P~vR?�u�hf�/gw�>��6��e��i,y����O$�����?�6��Hx���7�۵�ՇYf�(;�Ʊkrb	��3І=��Ё���
�1�f�s�N�+y9nͬ=��jTTEh9gNs�:��Y�>��n /�rQ�`��ͺ�86Q�m�O��F(��,�abS֑��W����Z�2;�@�M��B�oL��WP�s���HkH��Ԙ/��]�;�)F��DA��w���ς4�R����>J���8I%vU�\��tY^���������T6=:@�貊<��ޤoD
�Q梲����=��\������Xw�n��yb��{��[S��X	��<Z.�-Uk
��h!�4Zχ3y�Fo��q�㎠G�[3�#���+m����r��g���5)��eu[���׍�O�{��˄��ǭk�H$N����=�h���SA�p���x,,���'�;�S��o�mIɕ8� ����^��I"*�
~�#��`�7�K(���Y�*AD���sީ:����B�Z0�K����~w�~w�� Ф2��{g;N���i>�g`Mm��d�~�������W�޹K��2n�Qb3<����687��v!�Ȋ�nǤ��(����@�W`ʸ6���ŕjl3��U�����W���q�*(+z�C���^�I)1��iQ�,��9S�����7����?�6�iJ�L&���l.���J ��IjB]��Õ��,�0q�4�ĭ�3�.-��������ae
DX���$�-ޔ����^��&���Bsu?�Wʦ˂�a�ll��Z��vL�i����}��J|,���?,;UA��DW���^%E/���/ l [Z(��h~d�=7��1�zN;%���u^KR����>�;d&�S�UVi-���xlJBW��S.�1��NUR�s��9�'Z�C�F���$��O��M�$��V!�jeEH��9��VHܲ�%E���[2�nR�ʈ�w��	@4b�����a�>�n�hY1�$y[�>�����V��$�!�$QBv�2�2A�rkT	�!	��Zx�v��W��W�f٤{O��l�,��������M{�X��z��T=������f,�}��Vc�/]Tb���	"��O6.���nv�4v�93��m�H����O;�7(MBR�u��?2҆+�w9��`���x��T����z���n�bk��m���}����v��`�}km�+�HP��ڵ��mbW,�ųQK����VΤdطC�~�1�й�z�u��2��#u|p��c�E
�L�9@磝_m��!2씵�s�7ǒŋWA���n�qw#��,x?����t�N�}�TF�pi������A��U��ʳ�74s��g��o�	R�D��R��]+
�3�}v�vG�.�KRTl���D�:77{��)�w�<~��j]Z.Ҋݚ0�t���^�^�"zd����	�������k��F0UdY1Ɇ~�>���p�|�b���R�goRv�R��R�h^$˗2��6�ȳ��RQ�س2�L�0�_��l�*��|tW��E#�S�ÞX�:����#�!ǆF��Vwl��&��[��uqd�x��kU�Rk�m��1�W`�ˊ��eww�E${`&隧/��	+zm��${Qa��A��qTζ�߿��Д9��*9����'gH�_��@���>����"Tb��E �U��܇�J������#M���D�3f�3$�y):�O�qh"F�lo�5�(�� �{wD�PK;q��7fN�@{���h��첏ަx�TO�&�So�;��_�����[�L&aP_ҰP$���{��p�E�fr<Eg�x�VT���]l��D�����V�z4;��pi�bѲO������dβ^�w��{�hrm�(e˧^�ٻ�r���B�7S�~Is�I�fό����{oH�ʵ0[���?4(y Z�b~��m].ت*�"|�����C74]��Sf�ZB��Ѡ��j���w�7Hϑ�`	���=�7���e�
*-�H�l�l�P��}|��|��ݽ�c4w���]�e�e��3V	�S�d��������������U�gz�w�o����S�ߕ�C"��?m_~�F(3FlF�9��{��Bf#��� 7�_D]]�km�/N� ��G�����5Kn$�M??X��,m�h���ǆ�#LQ�T"��$2u%��W��E�¼3;��%���O�>�}�]��Q��k��rU�w�~�ݿԠ#�Cm�&�΀�gb�B�N�ޤ;�����
����+9��)�T]:��pt?	E�q؈?]l؋?�!��y�/ߛ0TT�c/���^9
�����R�5�n�ry1Mcǩr�z~,>��u�(7@���.���>>�.�>dﻁ�s�A��ό������;GN7�I���x���(����f�0|�Z����6��tP�d+�9��޼��`1"���_t�[���	N��-�a�ￗ�?*��i!At7< �_���C��"#����6�(��Ձa�o��,K�#�b�_� �s�P���&^ V���� J�R�8�?.��n_�D�
D���h[����{�W���[���h�J�*��Կ��9x��P>��-\��rMΨg�,�~�g�$^YG�@���4d�(�g:�@��O2���8S� ߳���ë��9]�L�=��C�Ps�>%#���w�h�VV�$��p���ҏ���ύ�����[:E�g�A��qf�f���}���ݧB��� b�@t��;2�b����m�'���e��Vf����C/e�S<���B�p��`����'�ϋT]����i�y���+J��X=�:1�������6LG�?+��ڗ7���p�QL=�|�-�6~�Sa�}����?h��qh,[���T�S�QW���Pg��|~�'�ʣ�J�������q�M�I�c����L/�]y��������ǣ�K�ZxIk���'/�����'�g������ߔX_��&Z�Mkwu�i9�;s�JMG�K��3�{}&�EcZ�˃��	󗲏��v=Z?X3���x�7�o	B~����d����fvK�o�*���n[��R����29�4����df6�hl���r�14����	����'�(�L�sm��:�&�l��it������k����v�W.�|�,1:@�y󻚊�[hY/ð:}�k�m�ua�r�ע�\Ӽ�O,]xb>KM�͸ߘ>�qg��4��aW�;S��nq����ܾ��6��D�H�Tu��F�*�_��sA|��N�o�.��.�!!��;��LrI��� ���q�B��ɺ ���<u�D��<ǘ����"_
~`�>�'"H˭c�e�$G�W�0)�Ȭ�������<Öz�u�����Cu3мΰ1�Ÿn��5���笍���Ź�h���w�\s<�v��C���_(�]1!3�U����nv���=~�����b,EU�
�cDg�
cIP��"���<�Z�Yu����½JN*7���|�$�Pr��1N�����\, ���^������4X�ZO[k\7~����cT��|��{n"4�v�I�'�'�����ĉpn0e��y���XP����x>��Q���qi�/Ђ����d�Uv��k!�_I�kj�?���)xH7_¹S\ëU��`��\�p����#/�Eg��n1X��3�e�ck��ԉ��f�gic6��.ٟ2݉�����]����7�(k+���S�l�fΐ��f���s�N����	gh.�c��޸h/�B��v�s��WBw|ǾU���Sx�h,%j�^��~g��Ժ�`ڃaRlͅ2��;D}p��������ɡ���>��.�,F�v�)�K�i�b�%|��Q�2e�f��	�z���1�������r�DO�@��.Ɲ�Q�/����⿭	��}x��nni���lY�*N�	����]4�pt.e��3�/!���(V/��n:�R��X����1�K�����#����B,G��d�`MP����4CO�E��C�
����J�6D��&�{7�������pc���4v�(%���+�Ldx
��^	f��,V&�^�{ɸ����ע+'8.�f�ܤ;K �~�Wf�}�W�g/4�;KQ���[�RH� o����<�>��c��H���u����o�d߳C������N]A�P3#�D���'�A찌�������W����]����Pa=_hh4nf���I�`�Zh�ë�+������nC�>+�н�?U��C���N"c��JpZ�5u0�Ĉ�(�1���+�*Wxx�g�׽�A�Y�Ln���K��K�N�i����`��^rd,V��[%��ĕ	�串>��p���)8>5��~-��`�[��_(R!�!Y�G�j��.�
�������&lдzq�P�������H&�zЕ�l*��o�V���B�W��@����W? i�D�ME�A���*���9����T��U���u�ش<�B�	��'��hT���tV��%m�0w� U�� n�	�²��:lΰ6��}�>��Jc��P-�趁ƓPQ��j��24;<�쿁����Y�uN� �6�n2L|��c�Ze�������OyJ�I���u"�c�N�aϸ��W���
�,�(�Qe��9�_=�7�����X�	9��������r��w��o���R����)�ܥ@x�z���J̐uxn���>�&�«��_���Q���)�T_'�����,d��sDK>����zv�ܛ�n��s�!ӱ���V�Pgr�����b���\1u���*������E)�A������ȹ�öZ�v�
�wc~�����x�jpY����G��]Y��5ٓ���=�dӒ��#A�_�gWʻ����p�\�=�~��[�B��xZ_#��\;�局T� 𭀓�mr����;��"w3Ȇ�&����G�{�Κ��vS6�=��!�D4�uY��8ס�/8
�Bk�ˀ�"i�C�e}��M1z73A|Mf��ҰY�z�@y��nc��~�¶� �ڟe�o��<s�|Cs*����r���"�۷^tS����3����&
��P�p��DHA�yj�'��W�َ�/��
R#S�F�t��b�MP�L�Ȭ����?�ݑM�%�>��B�-�����~�:��Y��CFݺ�'�FH��m/���&]�cK w�4L�������c ��:��� ����ox��� �c�l!#�}��χ{�<5YPk���
�&tU�������.*�O��*���0�����G2M��IPd���H��@g
�BJ�'V������d.��o$��=�V�H�{��9��--~���5��p�s<��OA��	�%=7�T����T�Q�v}v̄`"����i����.z�����UiJ�w��(«���q��� �a��]�*#+�Q-��Q���uZ��� m{�ؐ߉qة�i�������:(�*x�j�b�|&��;�_b �����豙9�R�����qx�a;a�추}����s=�{����x���4>��&�G�I����(t���v��$���?�J<A{춤�7��7��YH{��.HQ��y���O��_��قt�������6��%D���1��'E�	���]�
S���܃߹��?�Ci>4W�Cw���rg^��xڣ�v3P�*��LD3����������{>S�Z�ڙnX]��xb��s��Q�V�R	���a)�-�[y\����B��뒔�^��i�ِ=H��PX�
֣���/�|y�L0��#�h�ɁkWf��<�Fח(��SRj%�|�yø6��w���hc��=7����Z�Z��/���.|����Ԃp�-mݝ���:0=I (��D���5�Ѝ���#�Z&~x��_��)��`p`��&(Niݧ����w4��ܲ�o=��9�����TBͧ��o��_�� �Ss>�Z)&�+�Q��f@��VN|��i�a�D���w�A�~*�-%���f�q��] �㷂�uSw��2�ED�+���Rv4#���y�VD����s �`wu��Ai��ϱ�x�8^Tkx�B��&�=rө6Y�hH�P�F�YG�U�$�Z)����ۍ�.��gO����.��ʼϠ�5�7�͖2R�����k����n����?���T��=��h[]@�ր<68<5�y0���H}�a�ƿ6ȱf�����z���_����y�\c� ��:(�2r���/$�Vx0#���Y��ꚴȹ��� �:��q��\%,�|*%��.�_�S"5�����1�K�f����� ab�z�U�w|*�� �G8�u>+�?G�]�Х6H�)��/$H��hOp��tZT��Xj��Q�OQ�rȭ����z�~ss�|E&YF�m��}�R@)�3`�+��F��C���@�A���x�J������o��؉q��5��U�.A�,���O�8�����kL����u��tR�f�C�9�K����Y5Q��f��L�kf��%��,HF���'j?��(�+����JI{�����A^̪�:����>��'�E���Բ�SÉK�s������0���H�6ۏ7�/����=�~W*{�>�B�;z*�?5��zq�v���$UR����BZ�d*�S�(�E;���=�OL�`^�ߧ'%��A|[�V��‶��O�/��������>>h|�s�]3w�i�o�\9:m�&y*g�TПL��ܠа�4�M�v��&��lt�;��XP��f�a�j������t���X�r|$_�XR�3��y�A	~�k��I�˚��g�g0}���ᆪ>�ϝf��#��h���1�4�[9��.�,���c.q=�cQiD�"�:pݹ�Sr��u�6�3���n pD��DE��8)6rt����'�p5N���ظWt��ҹw�?A�6��ā=-�#��V[�>1Y��q�󠎼�Â����B�u����v�-�3��
I�r�Ӯ��[��*��F��#���@�~�x�P��R�/T�d�����10�=?�� �R�ٓ����I96.-271qH�.�vJ`·v&?��{�s2�����ʘ;XW��JR
���L�Qv1�>~8�B��\�9Z�38�Q 662��6����(.�c�\�|wV��y-��1n��8���G�e*��}b E�u}�������eϞ(�L�Cς�&�!��V�Д�tg�n���lĳ���,�EJ�YJ��v��J.���v�ƒzD�����P�q��<�w�|I$28gBf�o m�[���פ]f�P��l��ar�n�ׯ��-���ySnG������M�y5Z�xGZ]-�dP
<s��a��B������tZ�ݙ�w��x;�G��T;�R�`�dW�˧�ܮU�O�8T��i6���ߕ�)R���E��(ʺ�&�>����o�
��A̭�X%� �uϩ�<�)�Y���a��U��L
��a�:l7Q��Ɂ�y0���T�n�0E�����\����t#������k܏7��k'��K�j.ж����?�Q��E,�B}H����&���� 7!�C���ă���]��Etg���7;�)d�ڠ�"�K~I����E	���.C�l��,��@���;�����&����K�8�]Μ39�� ���~T��?��mOj*��hYMڴ��Z����(5���ff�i���7�߱���F���e�ܷ�;>1�����\5c+�_���l��eh�4-^�O�#��R;��MM��,��8_�HߺN���!`���8j��T��N�$��� ���WAk�Y�5�H4�M�u��Ű���������Kdlԁ��R���|-i��p	����4�x�q���O+��s��Ccq�،z8��T��h��3FpP��l-Rk`bbҎ_�VϢ9���~�ف*j�h]@��i�M�����j}3i��.�L�⍸ۆʒ��g���?R����
5�F��SŴS��G��&s�%�؍��[=jHڅׂ�f�%��`��:�V�(V�"8T�s�MA#l"�X谵f�hE�W�q��*`P3Y�:vtkr����x���RvxL��������Me[�����+�s�+2
�� ""J1b(�0#�:��A��Z0�6�U�Q�9�HW1 "E�^"�`��[B@HI�PB�w�s�}�?��|���|��>k���w���0�E ��b�>���f�}�J׌Ω혢H�����"�(�=;)�B�OG��h���[�ƾLÕ�[�i�e�6��!Ơ��LX'R�����L��*���#[ ���(i�@�M�Ǔ�lI����w����*It�2���_,�_qi�������w��_˪�峁˼(�+G|4G���>�5ޠ�Z�k�뎩��ʾA�6�IO��K� ���i�چh�S#1IJG��$�3����x��;�3�f�~�;�H��o�鿁3Lr����a;'�Ľ��X/tLU�:����N���+��A<����N��j�Hc"?jo��\[d	��mp��F12<0�67q"�b�%�)y���|�&���
l�ܨ=�լAY�B��M���M�Lg�OR�tZBC�5�W_��~B<�;�ݝ���oz�����z����K��i�m`��k��ȇhّ����� �a^h§��U��g��g{����7��������vz�ޚ'|��� a"�g���`����SV�L4�Z�b;��]�m�c	(T��г��l&L͛Z��V��݃ڪ��Y���zk}��+-��L�Qj�`��Us�����=4i*�ܴk�L�U�;��HC�Q�x�4Ӹ�O�<��w��ʑ%hr���HΛM̮�>% �䛚����Ԫ��	k�k#�3Ea���O��{q�~;�Q�0�-�J/V#{u�����K�}:�+�%vh���L_e����f���;n�(�3�f�F��W�����������Zx�BWؕ���f�of�q���Ӓ�I�v/n��[%՜/�ܨU4x���R���2�gO�.�G�R�p�ގ�q��)�6 �kY����$٣��#�/b˴_�k���c�������_����HTF��F�<cN�i	��e��� &r1�Cqdۼ�5n���J���7��ՠv�k]+4�_�q�ablxX"��Z�Y�m��uL�&1y��^�r<��Uk<NtZX@��e7������ͨ`�V'����˦ui'�xy}c�s.D�#.�@��U/�g��h�$c+ҋH wt;�2�n��U6� ����|���z���楳"i���3_U�a��ZV��\�Ò��K� ����v7jxdg����L��5�@�F��U�p/Y����ƍ�S�x�4���y�7�1�}�;�7�c�t��o�ε&Id��vSb����;�ƀy����x����ܐ��dgb�a����2Ȋ�[3%��W�v*�x��-�(����o'oC�ܷf��M��N���!�ԥ�YX��")��f�w�:�e���r�pc5�#�a��������u��8R^0lQ��ޮ����>8)H5T)G7m�
5�o����3y�aQk3c���#��&�gw5*�3a��S�޾���Uʈ�a��S6;�[��ns�@U�Bgc�����EbXf�� ���jO��[|%ju{Be�W >P��p�V�G�[;/s����*)]o�>������aL[y�
����{���4�s$AK����c���g*���Ab����TI3�$���$v���.���x�Ǉq����j�"�X�&;�Z���1��=�`7}k���p�P%�=<�ȕ�{�Rn4��|L�$���gMX���h�`(P?����-���G2�{iG��R�?���/��쎥���4�z�_��~(a�%%xCh�`MIG�,�7���B��.�"^s��h�w/�[��4�e�~s�Ɩ"�>�5p���7����kヮ];A�IF��!�`��3�񺒭dT�F'Y�2>����SV��Ǐ�ێ�t+�R#�k˛ƍI�����7�xc5*(���|����ONĊ2%��%��ȿ���K�c���e�SY���rT���\�U������V����"�[_�FӱZKY�g:qhs�+P8�G�
����Qb0�5dP���2�C��Q�z����&���|�ٶ�~s��iw-Xd.���Cp�B��k�y��Wg�z����A����T��3��+F0<��E���3�=�=�"U���� �(6����d��g�>5E���t\� m���;2v���"@* ���I�1��4�	��U�?�Y�˨�G�����*@���a��%*�O!��v�U(`I� і7kh���v�T:�ٖ�g�u|k���l�\,�3c&��x[Hh+_Ur��|������������H�L?#�3�5����mc=
�o�!{���Y3�/*�GN�l���	.��=|aKC�5O�kd#]~��6h������NjD ,-F[}ܪ=*�V�I�A�Y~�]�ۡ��6Ho�@)ϊJ�e#ms����w��є�̖�ϽiM~u_�7�Q�f�C�s
Bd�G�J��̳�1 g�q�wO��湠���_}��6�\�ffY����ؾ��h�/�Xgě����E��,]ZPp�-�@�� BmF>�%c$�j����ѵ_h��dC( �}���v�(g<]��K@<HZC�]뫵uTmP��NI0#V��D�5����7�ۊLTȝ[$��ɜǀ��
iO��%�^� ��oղ�0������.��h�%�'�g�Ɗ� i���~�Y�!�k���7;��� 
 ����Av�c��
�8���N��ϺcE:���ϻ���1ό[I�K���:#i,����My��p�v���2T�Yß��o)1	A��aF�������x<�q��(kU�7D�V	� �M��:��D�^w#�0(r���O�,���j@�
��0+�����
 |��i���p��f�-�E��J��Mɍ��K0j���C��~f<csb~,��xDŤw��1%gp����gd��c���y��]P�2tg|��b���ț�� Y�S��8�<i��M�(��]��x���.� �ŌO\�w:��AO�� �?���h�2�c��w�wu�H�W��3�Tέ��{�] n���rݿ�a	�O��*�~i����|9�>B�#�La�z>>Hr�!�q�oܛj	4|�|����sv�d���#�������J�@́�����;ekm��2@Bu<FK��.إs!��E3����@~3v�~��A%�0@�G��#n�(4�k1H�*�W�Q'@G�yP,&�ghj��3 �W'y,���2����Qa�MĻ^�ѕ�d�F�����2��a0H���#�Z���}w��Q�ڋ�i���e��n����p��砀R[twl�O�xf�մ151������/����e���6��d��,��T�>,Z����{A�}�?o7L4�S����� ��u���Vgu�����z)񹒳#�
��$��Ǩ�mFM��ۨT3��1��o���r*B`�ǩ��l�9� ��!O����b[=�\;�(&v2݉^)�-</�"�e1�E\(��}����S�&O���E��)�\��m�B�  ac�u�bC����7`��Lb�)\�=#ǣ��81\W������� 3:f�Z^9�cw�[���� ������6,'8��+-��r��
��pQ>**�����
7��,�+�kw�w*/��G�K�` ��"O�Z�zP�$	cq��V���x��d`
�]����]Rfa��LE!Pt=x����Z�/��s��-CI�
n$$�B�� �h,ù>n�u���z�ºJ���	 �v"�!�~6LU��^�͊�%��Z��K_ *T=��b$/x0�0�?�>Kќ����B �M'�T`H����j�SnL��8Hl3_�>�m��7��t
;�a�AdK��}��&�z���C����r��n�Ҝ��{q$��9� �+���\|�
c��ٗ���`�^mG���<ި��"z���Y����N�%�\����>���o�!��?�pZ7�`�ô��wJjn���ܻ�9�UL�X�R��YR�_��:���Pٖ|y ��t}�i������F�xC�����q�'�C�Ca���5|�O��Z ;K<Q9^(1�����T��W��y� +3�e���t���!�1n<�W��Lu��v�!zwl˨���2�����Wq�z��F���3ޙ�� �s�,$f���+ ��(��oj����y�W�	�.��Y���#xw�Q����1�  O�C�;u��tl�(�󭻘�9�co��e�j�T��y��1�	zH5#,��ɡ0�IF|�s�͖�ɗQ^�����r���n��@����o0�j/Rf���;Zb��l�c�|vm�tc`�P\/Ā��]� ��!Ts�\�'A1�� �(�x�S�� n�ѓ�1�?�5�0z/叝�����|���a�X���d����L��f|c�z���8}��������3�ȗ0xL3^�"�m�$�c9F�=�<2
^��5D�eay�I١-�t|M���v���q�Co�z���շ_}�������_��_����o�Ҿ��+G������F���]Z�>5䁕�����__���չ&iԯ}`=O0
��J�7�w>v��|U~�0��P%�g{F�Os�xGK�D������ݮIQst�=�]lί,?�28�e�ш�F�O�v_,<�-N:�̰"5���[��^m����C��aO�۶�a���N���A�5T9rW�-϶���}�6z�®X\ά_�x�Q@uqĽ;����9����E~�3v�J�OB&�� BnYYF�h�R��r�|z	�E@��_g�i��-#?R~p�O��M��o���Z�0��@�ь� F]�	�����6��%$����~0��O��Ԩg��*��{)�1��3UF-u���»:��L��	j�iIl���~�HI�����v��K��� � <����u�L{8��W0��q>�	��a��!�'�D�#҂*��@�,O�v���9��z ?F���e�'V�
��p]֯�?G��,�\���������ǹ�'0��a�q��6�������x%0o)ݺ4��S��t�M2o)���=T�O��G�+��zĸ'˳ꍨ!!e�0�cN���Ӿ���*�J���)#�-bu�ܢ԰���O�\���T8�ed����h'c��i�>��v&��;�T�j�+�k^�����[C?�%F�/eK� C�tU�w�BdBY~����+���4�YC25~^s1�
_�T��i��1ة �efh�?9OO��z�u�%��|�?��nO8��"�ax��.U1��y#YG�ͱ�������R��XF�G/T��H�ϕ��~;�~�$�1�iL�Yܕ�u�X@�g���ZUG��eU'M��? go�o?8��t+v��E�@b���(j��ä�'�.�<Nh����3��gB]���	=�>���}���U�Y�U2������|�)����^4���{��Vo����VVgq�FvD�t��O�:�T`*�&X�G��ʱr��0��LO;U�>I k�Xl��ʕ� ���]pWb���$�ID���Iv�i�h7�C7�U�"�p6�q�w�U�S��Y��F7~�"g���4�rgUݵ1��%j����C��1�y�����9������39��@z�b���|4�Ǘ>��er�G7~��� -���<��q�9|P�kݎ��Oһ�:�{�ʮ���#���B�V��3��/SaǈbdiA�)1z�B�&ܔ��V�6�{��o�d'*���F�&�7b:0�ڦ���akW����F*<�ꋿp�j����6l��ZL����(_�3$�ߩpZ��q,?hߓ��KH^o4\��IY�n�$Ͽ�ɃG�0r ��8+ݎ��uv�?�+��o�h�\�R �_K#�N�-7���"�^��k��L鉹����e��>VР�0g���Y~�)7ZJ`�
��<K�|(����Ȗ��퓻�\�b��d$��ػ��s�m������1h� �T3�F��y��k2�,m䫹ſ8c��r�ȷ���i\��j7 Օ$���n��B�D�[0�s'oIVC�IDH���
���7n�į�ni���շА�K\Bn�E���Z���b"�8����[���[�A�/	�V��;`�U�������ḱt����'Y�b�\w�f(����1m�i&��ލ�(����!�dH몥�[~��	��[C0�*Վ��A��pȚ{7j�<x:��(HHu4'�[fP�~Lz���P0v@;"�2��G�4ǽ��цG-�~�j��F�z���.�ye%�]%�_D-�F�7_�ʸE��d̶j6]�@2*�O{lh��y�\�N�ҝ��R7Z��ep���xu��(�t��e54���@�UK�2A��1����]�	�y���o�^�*��D����9	F�Wj�Ѩ����W���Q�D��T�	��	��8)W� ���;�6�6�
0r��lK��s l�ү���`�x�Mo+��,;��,�ӊ���w��)��]��F|��]�g9�C�+k�J�8�B�jA�Va(c�^`t��>9�5'
(9_}R�|2z�tX�o�Nk�- ����ֽ��{ҧl �`u����ͬۡ.G�^�eȻ�6W����O���7Q .qK��Qi���e���b1�Ϊ�㣖A���������k��I�G��R�I��f�>�l䀉/b[�cG���b�C��O�����}c�]��B�����1y�BW��4��a��~�6';���տ�V%��EMk������pR מ��4�F}�q�v��������/]m|9��55��YD2͎��$IF��������2�Y�VB������n+�%�ro4̑2����)}u%B�"�`���a�P�����mkX�Aއ2�:o}�������@������6e�ŧ�ڻjX��Q��v��ZH�l鮗|'�Y���)79��5|�~RN�%�7����e��Q4���eTȁ�n��F)9��h���!{��^�i>��FE��&w���G���mW�u����R���қ�U�6�v̐�����7Fv cO��M�H&��+c�fA�#���~�J��T���P��ڌ��Q�<�i��1�L
?�u��A�(%��^_����$�q�z���[��&�c�`"�e{�=dp�a
"WZ���z �[H�ߞ=�O��ظN�\v?>��d��<�٩ۏ���#��N�;� �P�:�H!D{�$�Y�HT8JO���	�8�j04�Le^��E�J�<X�c�R�$���޳y5� e�sh�����you;�|��'nr+����;���q�9䭪�<��1��Z�9��a� ��>i��#\�˔��`DR3��&977j@tҫ�k#�*��fk�ֳ�s�_�Go|٫$-h\LwT�	p�yX�{By���v�M��BVw�.�k�� �������_��y=4������u���%������ߊ@�H<^5(�o�2�0��՞�)�ҋa]Y�j�u �&َ����$$�4�Ƨ��[�0	��_&��`hq�xr�M#�z���uO�(��2>=W���U��J����^�<�>B�N`�aV�����W}ѻ]n$4�GG�|.l|��8�s?f���럚eT���SO(US�,Oc����2�FƁ��@��0(��d�ضn���v���u+��B;Y�XQ��	���_��!�!������g� �)����7��<�W���P�h��(�4�<ډ��hz�F7���=�D��eKRӄ�.^&�C��򋻋N��`��矚Qg��*'���׌�1�%��*-�Z�ږ��J��'9���-�1���v���:P֨�:XY�=@CXS�xC4��d�}���1� Ð�����+ulA�Y��J��hEQ2AZYv���l�Id�䞨jF�+ǻ�!#�~)� �ƛ�<M��zK"#�X�2ΠM�t���@�ȣ�Bj*3 ͜�(��p��a�2B_�R\]j�;p&����䟠8r��1MU�?�p��m�dB��)�G0�rn��ܖ��C���C���č�v>9;���v���(�~����٪V9*vE'�D�Q��z ׁ@/4x�B�[���ض��q�@h A����{�Te'Nv�Y5�jΧw�T�A$�q��0��(ޮ�%�3�����+'���b�;n~=�q��$�Ӓ�o�v�[X;rs����E,�Ez,Y��5n����_�|�9J�܄�L��KI�ƍ��HWn�o�U��+��r<���2,!��W:��?�~�d���d�_�jF#��C�� ��B�L�cY�,h�H�������Sɘ�paK9��J�t0��Q,O����]�B����T�|�AېQ�����Sc�)&�:(�{��M��3�!�1*Ȇ�!Z�=�hD��L��gO:���X9[�kS>�Z��XZe>�l�q�l������fR
I_��Q�,N�ș�}y�h4�27>���r�Ʃ|�i�!�Uw�o
jY�@� ��,&��+J>�{)�k�j��xH��Z�ԆN�ذ=�n��!1��˛�Ι؇WJ���ُtw�_qn~�*8X^R�='OXk�0R��>��9���L5��gr�m��d��qzϩS���5Z6�_H���Ĳ�S짙�Tu�z������`BV5�}�tsD�\���Ǩ��o�+�ygl��*�+'#���x�Ǭ��{�|zW��B�ܵ�/3��No\��8�m�\��j5cD1�����f��8y��GhPE��SǗ�Aɘ�~B��͵D��B� ��޴,� 5$&��Q�����֩Ҫ�R����/'@:T�)@N�sc��Z�Sc��-���d-�𙇘0s���c�6ɼ�WS�ސ�÷��Jaȩ�"4�����~�iT������2�G�8W��}�6\�n��}���������r�����t5�Yn���6�F����V�e�VR����`��fRh:�F���1�dxEԓ�f$3yp?kN�n���@SJs�<o���@�����u ٹd��[��WԻ�Q���T�a�P�N1:�u:��t(BT�~gkO�#~����&�2:�XF��Z�Q�����s�o<qaV��#�[�{XtT�<o]��p����⩛x�'���m��<�V�C4��e
)� Ħ��h?=���K��@�$��V��]!�������W���|(@^aR@x>�����%��񫔍�����(����{Y�AW��c��@�	�7 � ���]�a2в����k��-�N�a;����T�5'o�=�9�b�f;�קE%6Fp-��$��]��^O�=kQbֿ�S�������!F�Mû?�Q}���|*���⳨��oW^�(���I�_�w�����V��OƊ����v!�ш���U�9��n+�?���õh�vj�(��=��O_em���Gj�c��/�����܊�(5�zܨ�(�����9/A
�+&�~��w����jK��B-X��Nc��:�W��?�~��"B񄳀db.yi!��coՄ�)@�bp�ċ��ikM��&`9�
�g�͑{J^�'����GG�b+b�w��b���~?�(�E�MY���͓�lm��,������������g�n��NG����^f\���<�#��'��/���J}����礶��+��
�D�,��;qP��rُ�K��'��q�f���	�����ۭ�h�,�Tk;(J�1_��>��U�:n��K���HnH�ZIn�<y�Q Ej�(\F�_�cm��x!����1H�}�n�l�w�7\��n��;��&g������C��8-�[/R�����c\-�p�>��VW�ۡ�[)�hۙ5"�<��JRc}<�R%�B�Pb�~_I��l�Ju 7���LB��4����R�#��T��<f0(I�j�z+��Oj�)�Sm\&������ 9�a;l�H��a�h"�h�l6A�1�$�G¥h�C'�Zw�1J�/Ny�^fZ�es����Wݿ{w�Ġd^��9���ݠ2(á�����;f���Z��C���D����������a%���_M6���%�}��`ղ� *��4�ί7^Q�)j�2� &C.w9���t�F_���J�:��
����k�����bEcs^B�v
5�{<��t�mii��z���?�{�+)nF�7�o�m|T�m���^�𵝴�0�XcZnbe��Q����+D1�AMh	%�
k1���{�˨Tz���rg��<�I<*��)���*g7~�x���<L*���Z�+۔�ڤfU��vSӑ"D1iŊ��;m�3~�W�ӛ!F��~�_��}�\��j=�D����{ݪh,C��蟋]�"xx��}^��#�,�?̵GCNiI��q9QF���uy	]�i��P/55q�O���}�h^U�HXr����c;y�Ս	�4�8�Sw$a>ۂ�ɻ�b@�����?�7'3���AԴ��oǊ����r�Q3>dQ���F����T������lȘ#*z��'� +�J����y���7M�0����-�X9rĠEO�+7����$�����DE'C\ifb4�բG4�w�=}nϕB���>Մ�����^�C��[9�!943
/D�6����r�$����2c"uk�6�<}fv��	
��jX"։�Z{�=lH�9/7 �|H�E�UA��U\��� UjÃW�Ki?n��P��Z�����+f��ԆxN�K����	x/2E,���|��̉�v�о�,v��6+}Fj���4�]t�s�{u�Ǝ8�+�r��`���N4�k���(4}<~=���5k�}f20tjǓ��q�]���c�dyD�N��;r��/M�L0�}?(!`>��1j?�
̉!8/�G�p:˝o��v��U�A?�3"��x�!�(�)�ۊֶ"� ��[�0eg�_���-���R9,�"p�X� ®��͍���y����oW��؏Yڲ��?��+�5���@���;��l{�R�y���8���,@��0��@B�;-��_��b(��J�'������;�����J/�ڔ�#ϻ]�}��b�͛6������~� v���Tҗv�':/ X��֭l����;��n�1P����>PX��UMj�%lK%�%��.@�H����"ۜoDxF=��a/�
����tNT9�ݺI�E�?�t[��aɬ���R.Ʊ8��s}}���k.�>`���>wdW/��M��H�̹��V㎅�4��
	�,��Qv>j�M/������e�����ix%��uy���ǎW锂
ĸN�CD��R����{�O�P��H7=/7���O>���&�֨�+*
��{�4��iQo��b9@�4'��Z|�4{�H��iv�������A�n����>i�v�Q�y��({0��t�3B`����A��x�	�G�8��N,�$ �@Zb�!F<X^�O%���ԍ̄\�>X�����W��ʬݼ���L�u�g~k�|��3�
�S1s@h�\2?����)���cU:�^yy��lA���dV�kj��<zs����x�I���,#�@'�(�f�hF����L���p�79E��k���@���?��lF��d�z�a7^�5�F�fB�n�I+R��ҭWn����z���hi�F ����
�?�D��~.�g=����}n�ԅ�fۮ�
��)�EkN�Wo:��آ��o��ȑ���Xh?�U N�XӬ,O6c�=>�&b��,=W���{�T��#E��:��5���˰�&*�jxP��:0�g��%��2�ޗ�S3"̰�\�|���#I@m�)�;F(��83#�b��Z�-�G7aLF�XV:���)��v�ތL[�<D�c7���^����<{-�-�{����S���Ճ�@�I��sxfƘP�
�2KHmf�&u2;��)C_��-���#ݶu�o��?��Kvy�=(>Ɠ�-u 傕�]Ξr�3o4��]�hL?�n�ퟕaP?�{5�Y}�9�߲v#��/����g�٫�qO��E�x%�_Ց�����B�]Uv�����t������;3|*ŏ�樑�G��9d�O/�_��ͭ_��=�LBdd�Z�k'��9�լ�\�9�ň��w@���r�c
̙����+U����IFw��K�v�v^�����
v��5t���/~p��_j\I�75���&����`�D����2:����\8� �u8M5�nB��Ix8|�Y���P�I���ثw�d�E��E:l���Ϸ^�P^�h��φl>A�[ ˛O
Pc���0�������Wڑd[���^�ɨY�K1\�����0�Hm_;*�=��Ԉ���U�v��OO��
G��ː^9�̐\w�ۮv��y�NUp&�A����Qu���Ʒ��������UB�lK�u���#=`�#4���95��e8�|3~'v'5�x_�|)� qUv}��^��qQ/��#�je��g��ވ�@����bJ�5b_�-�FS'���3$v"Gr�nq��ה�R�����xL�*!8'��v���^��A(��'M�"y�\C�k��"��RVc�,5�x��4X�[W�^�q~j�� :�=(�nG���>ܴuu�z���l!y�lH���Gi��_ /R��*���'���uU�%�4P1��T%Tu �m���Y��73&i������<��)R�2Q>[ֲ?�W�坨��4�G�S�芖8�[ci�7�=}g�</O�Y�;7�u��U��q4�鲼���33�G������vo�8��Q}��$5|0�}�:!�G���>�lg�^<64c���A�m�)Y�	od�x�U(Tй���ѥ��䫒I�Ɗ����/w*�d(�U�~��K��>�K?)-8�Xj��P����9^���YyDsc,7GwEy�+Ɲ��9��\��� O!x�0�^�����D��@F����l�o���\�̃���6O0�F4i_:^%W��n�X�#��>9�~*SG"�XƸQ��ah�Ȅ�7G=�'7�L��9)��Ș�ЦM+G�E=��ba��Y&�mΧ��I�Lo��Z������iֻ��l�!�i:��{��$;�A��G��a�H�lMZ]	~Ӎ���bk.,%ͤ��/r>^��qܕ1�=�GW��|�B�u�n��#���zEmR%Z��B\(���rN�R�����ϗ5ͩ��_=��U�� �8�'m��h=������̫#�z���Db�D��8T rb���j�K����N?![?���b��Rh4�O?o�Tdq?�h��P(�V�ԍ����ʡ}�N�w�h0b!�>�DMG�����A2�Llc�iE�[tz׈��;��\����u���"�i<*��.j�����Բx�wV~��	���5K���x�BظG�yy�2ݨE:�'jST�H�ۃȖQ�鰶b՟o�P�,f5�:���>�n�Y���~+r]=S:����!���a���������T��F��3ٍ��g,��o*::�o�3b8�+�\�͈2���'!)嘒,op�b�	�Ǖ�O6 ������.g�Pm�*h��?~�4�y�hc׬2(T�|ҀUΗEkY-� 9���?�Ċ�[�(�1^m\ Hᮭ�cVS�oZ�~�`398�A��{�v��z�#']�8���'(a��Z�f�S�P�Tw��D/���t[��kǽ�ń4(�+4rH������j$�+UU�Zb���'m����m��)E�3_!�l&�s��=A������;��'�; $}�Z�����9C ����+�@qI�=�+u[�M�.���x�2�T�L�7�D�o������¨�^?mVW٫���(���I�$d��E�w#�k0�����Z����V�T��1?������Bڰۑ�]�!���;Z��n���������oj��+U��۠_���WPai=V=�kXDz�|��!��H��3!;�"�<�*����2H�J� ��o��w��P�~�oj�R"�֭� sj�ߧ4���?B$�?��L� Q�ո�Ο
HR�~�iu�˯^b8��S���$�+k�
43�.�6am|1�6��Dy�[�Am{�*�WF`�MT\ft1��J�!�{���	�q�i���O!K]P����4�<1Z� 	(%= ��"27�%�M�"%&�S��p������s�ܑ��1B1O-��KKTk9�~���Klc���LU!̧/Y�o�퍍�P�+��Q%#ϛ�NVU�\�pG��$4���v����r.m�f�Ԕ��[�KoO�7�U=�h��8��*J�����*�F#ga;>��x��^�Ч!1W�{'8xZ��J�g��l�tzg2�14R��(!6e*�٨w�����h����Uey�����j��3.�2GПԚ�3։/XVK'ͯZ��sٛ�l�f�k��,sE3��F����٠�|{��|�[�c��
�d��y<�pr���d.����x�|X��;��GΤ6F�v�p�,X<��l�A�5��/�/0���Yo�JWV
z��8n^�}�ǜ�ңۅ�!�z>��͸sT�y^]��j�"[2I3�䤦.Cd^��{*�lvȇ�A>�0'�=�L�>G$,�'VD����pԷ~�iT��-De�^uZ��}C�k�\��QG"͘��q�{S��5��O�h�D.s�*�n�,qI�u�&�9@�PIq���S'�l�^��`=͂�B(�Ca҂���=(?raOB�}�`��WH���Ygd�%K^��X=b�]�}�^��гzT�R��D7���M��+�O^��Z�-��h�D�uܝ�P��V��iY�� �}�e|l�U�5,����B�����$+�z��aί�I���k��{f�Y#�r�a����]��d2�$K�QR}�C���Ɯ$�ht'�g��8L�����b�J{�U����KDft=71쨵e�F�"���ԥ�{�)W-ԽS����-�P�ɼ7�Z0��XX,l�癬��}e�7��5_%��28[M�^1�H��@UU��i���2 ����21>��Ȉc����fh��)	{q̯��@�~���E�rZQ��^�Ȧ�}Y��*�v�4�����%���R�#-�I/�Q:��;�lS�n;}����%�k��W.{�c�7}?n�Z�;��'�q�N��#?�����5R��{~�~m�� k�I��[py�_�O��uK}���Qj�.t�ￗ�pZ�S���-���B��/��B��/��B��������oRRߒ� ���B������S�J��
1�.����ߌ��v���p�c�OJi���no����5Z���.5Գ(_<�>�V�xO3rc��`žK���酱��^���>��b��ӧR��㗖�II]�i1�zG�(R)��MMbo������B��/��B��nΉ
&�#K��=�I!ӛM���������Fj~~��y�*�P��V�pc��=�_d��vg��#�S���ۤj?������x�tU�[vm`�z�\�h�)^�9p������K�Z��2!y�I2�g�e%s��yL2�%ɜ/>����_|!���_|!����fCOwJ}��ڴ�e���k|+�f�z������x!c�t#������w֝mj|\�,�,��������K��PK   F�X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   F�X����H   C   /   images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngC �߉PNG

   IHDR   d   4   |l��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��|yx����=[2�=dOHB6H���Ȧ�
����R��jk{�t���zi۷������R�*b�V@TY!@����=��d��=�L&$di����I~�[���g��9Ϡ�Y�����b�x�Ǉ���'NwC�R�j.�s��u�B��Z�?q�'-jJj��c��c¡�v9�v�w,��G�O{5:L�	}xߋ�mgI34�o��RB��h-��%C����v��:as�q5��Q89O�2{{Z|؟����,{r��
�:6B�U������B̞1}�������N���*�Z��Mya�������\.}2��Á��V��P+ZL�o5M`�����3�)++3(o۾� ={�ɖ�j,tOrL�_�:��E�]�����������S�qy��Mʰ:7�-Σ	��my.�cA�	Ĭ��Q�Oar�e^�3<C��Y�e��w���k�5|���Pw-��X�'V翐�����mGOgZ�.��e����@�� B�@t�Q�֪eR6��f�賸au)}~\���e��^\���RM�����FNz2�:��i'���G���E+�AH �F�9D��59�X��5;e��DJ�V*����8~z�ɷ&'�{%8P�����V6w@�V*���j4t<5!6�ʖ^�4t�	Wx\HU� c�MN����H��BhH04�h��h�Z��׏��v�jơ�N�t�`�0|=0,�H�����c0(*�I�t@���p{!���1==�s�0-k<�b���@Q@���fC���ӭ�8^݂/��Q�a�٥5�"96�/k���7O�}s[��*��,�AV豿��������7�"�X[�������i!��T�wAI㓑7m*V,�A�ށ�GK�i%���p��Ac������D�.h�k�W�I����~�(��f�c�iț<������zss�`�utuu�HI����k���U���� �m���Q�D������*�
n��Wb�j�3�
��	hii��`�
!�������T���a���������CxsW��c��'�e�A�ų"`�*Fŧ�jZpOON�����W"V>/y�%!xx��#8�h)���D{{;��܌��^!:�����0aRRRI�187%%a��|��{��8��.�O��9��zΚ��-�I6���+������������ݻ�u�V�<yR�Ɏ�d�J�PZHFF�.]�U�V!++	I����k�?�8�����e�U�5Rg�w7Y�ƣ��	�"'#���?�>���
M&�yY�F�҅�����~I��r~pЌ#G�࣏>�W_}%��K��S	�������E��zsss1.:wݴy�����wa{�����I�ya0R¼x��B,_�� X�"�oߎW_}� 5�e��F=:G��Y,�8q���X�~=��<��Cb=�����"�����r�Pغ�f^��һ1))ڀK�C����}&|Yg@u�Opc#X��S7��{�,CHX�X;�?�	��n���3�*��+��y}�x���
Q�w�yG@�я~���Lg*��X$��ފGڅ���9���T<YƳ�Q��Y"q�������q�F�8�d�PrK� MVE���dF?i�iP����_��_�w���ϟ�I�&�?P��ڇ�]k�83g-2���Rf���$���g)�C.L�g�ñ�%y�B4�9ߣvS�䖟X���X)q�l6�7���/��Ʉ Zg�&�ؙ��
^/���t�J�`��[��o�>��7��ʕ+����_~�k�-��q6&�&�f���ibFSS~������iub��� L�LG�����F&Ǉ�h���@{[�O���|�V�Eyy9x����X�b2H{��ף�孨��H�c0��`4ۄy�"#)
��:8u�A+ٍ͋9�0c�x�t�CK|>6"�m��n��¼t4wP\݊�-2�G�����߂x�n�Y8��r��100�g�y���D��`�൦f�#�,��(��C`��Bz��q���vY�^�Ǐ�cqs=� b���Խˡ7��%6ӛ
�(f\+��������i30uz��G1�?%��9-@�]\,�f��T)�ع��� �F#�q����Ǵi����v<��ð�Ւf���z�"��ff�AO���!� ���us�VbޔT��eAv2��}�
'cJZJj�x`�l�,vܺx�\s��E��?�Q���o]���q��>��h7��C��&�!o�L�Q�~v��1�x ���D\�R���܂S�J`"p���{N�����GJ�<~�BԾ����HLF��G*��U� <"2;v/~0xL��M$���?�ȄU�O9����Y�/Qdm�������(!�_�BX���������n�K�Y�y�t2o/lD���l�l[��SR����퇫�EI
rRĪq�dQZa0�SSq����Z�;<XK�ha�9d^��5��ƙ4�	���� Afdgaz�,YӅT�����dM�QQ(:p]�bM,K&9�/F��<ܽ��o�aG|�y�z�Ǎ��fbJN���mۆM�6[��=u
M�-�����u ��i���iBPp%N��I#<����7^}�>�P��^HB(������=�P0W�jw���G���0g��N
�UL{�	�����ാs&���6��d塺@Y���:|t����Š�!�E����)QX4o�ģS�Nᥗ^b�H����s|5�`��
�u�'H�3���%2��x!����=��)S� �<����`��F�u��s�a@8�'�����>�'6,(�C�I���IS'K��+X�J�H۬V�\32�
$���<AC~ۋd���q;�|��K��c�	|7�p�fcav�QL�B};�,Y�6�-���pk5h�6�bs�����(�m��RJ�0�,�&�<��M[(����u�`�,C���f�x1��^{}}}$�-��ř��ȝn�:���!�ޡШ��{Y�V���B��OwJLe��Ĉ�����3SQ�I�0À���ɈFf��{׮]�Y[8�O�1]bSvO+�&8�%��vv��7�L>�4-��$��T,�����g���Ѽ6��P޲���֓� ���LEc��fsbDPf+9R�$����Ҙ���51|o߀e�^!I:̜�-��4~�Ν�r)S��|!*~ː�@8]kHl!�TС$r��x�?b\$&Q��x�����vYI�����{��c�Q}���B�<2����l��ux|�NԖՊ���\��`�X�� �W�J@#Ka��Қ3o.N/����~]]�$Ry�iH
/BC����$^�)J���tW94'���G�+Z׬�����?���az�������n��p�.X��;�e����jQ���Z	�LKANB�֛I�J l�Q:%rғ��B�؟2�<A~�
[�m�B�g���_�j����3y���db$��u��=zT ���AV\��p�5��C�ʃ܌DZ_ �/��R\1��#צ䎥�u1��3� �:>�aוH�My�S�$�˗/��w���}>�bB4�����\��:O��:�؂�'Iʔ��-�27���ޞ^�EF�ű��H21���Zy?+ ��MYc�WjpHP"5!F��K�O�<)w`e.���\�^��5)\^���K�Gme����Sl���'FQ���k��R�@}ȣ��U\	�I����Sc�p�e�����5(�
����v��V�K<A.Nr�NK~;n\���Tx�еJD���ߜk��b�j��Q��� W
�m���?}����}��a �{�A�/TK=����%�`���ݗ��QA���6��5�`.E(����X	t�@J��[׉����!-�r�w�}�af5�!����u��Ā��:8V���rrhw�`YBۆ�����-�@��O�Juق��:���pY��D����|_�0z� p9}�Kz��{����0 V
B,,h�����5ea-%��;i�<h|��XK�W�9�:����؛�{����8씧8�\���������/!��'��i�)��}���X9q1��N�P_�jw�)��Ff�qXOLL���o0צ���M�R��C��;)	�Sk~'�D�tW��p|%��D����c6L}�UV�v��a�U�*�4�r��^�N�db�M.ޚ-�=Oo�	z>��D��ϻMNt�(�NEzz:"�]q,��%ם8��=�)����b�F��Q¦PKi�=�շ����p�qM�,\��O6�=h�����ڒ(q�0V�F~���+>�
	̸��� ��2q����;?��w�."8��}p�)��B��Yݨi�cf�4����P6�EEF���q��#�&�G�'�����)��mX`���K��]�b���={�\�Mϭ�0�J��݃�is)P~�+Ic�����L���66 ��U��O%�����
�`W�J����A��FC*�{x����%��l�����cٲeؿ��.q.\ ~����,#-3�Cp�|��٘��.�x�:�a�:�;l�-s� ;;��@Em#�\���"�c�� &6Nji����F�]u8y	�q|��[Ɍ�uaP���rD��$���5��g���Ȁ�hjmC��$uAëf����Pd�p����E*��z=v~�V�^��d)D�R3ӥc&�+Ŷ��S���N>��gS���r
g����K��j1c��Z��\Y<�&V�6���:,��EAA�Ν+JȊT^r
�/
���J�Z��ű�<W9X�آ��J��bs��Sb�L�V�^����1v��
mnz�Y�E��6�����Id��3�>� ~��_I�ݻ{�⑛7��Cu����}Z#�`4�IBg�Х�D����<!+e��Ipsб`��N���{�;G5�.u\l�$nڦ�����;3O�G��?���Ue����c�C�x).(�P�������ix,�_�B+[���>�2��6l/��-QC���C��6��wO#3+w�y����U�-��$�͞�#����W��9Fh�>6�4�Y��Ox���C�슷�<���B���Al�u�F�9E�1�s=�� V�E�z��'۱�D��?Gv��{��K�PY�I!.ܐ��s"t.~��G^/ˢ��hnh����~&ۣ�7>���hTg��(��M��N6l;���(�췿���5������o���� �����~�Q�P=�'�A���ȧ)~�q�z֬Y"ރG����U4g��gh���k��i�F������T7wK�W��C���h7+�����JCTL,�|�I���ٳG@9q�X����dS��!~|p:QT���&���>�(n��f�7����]�{U���O� ��=Ԅ�̃X{�R��*6皚i��۵ՕU�6#_�V���=C�Tu�:�(^�46����@��׿���.�����K���::v�ă�CT��6�GZ�	Q����'���'�s��[��C� k�	ύ[�g��rf|�?�{�R���?����,�RGk�loGVN��Wt�[T@�(���O���N6=�e0�������\<����l�C��<��[������,B\T8
��A^^�~�mq/���İ�(���>��01��p�0P�����8@ԸG,�����yO[�ڵk��v=^ܰ���"�Q�F��I��w
{,r���zS'QgàPU7�E�E�D�t��}=s/2T�%��9<\�4�����<��|V��ؽX�l)�������f�͛7����?�*O�b%u�Q�E����k��$����o�y��`��!�¥eЄ�l܁��]R�:{��e�u��y����4�ysfc�ĉX�n� ��[o�����4�Y1BQFm��I�֬Y�'�xBr�yԞ_�16��WFvC\�	"vc���[G��99�������ơ��$J %%�|�ь� -��c��/�)��{_ɽ7^����b)LO�Cp��˙<����ԐG�[��pn�.�c�op��u?�+;��R��A�%��_�T�O��9�6�K
%���?�Nז-[�^__/%��2È�[/��-K���1�PQQ����������B�������;��/��~�_����za�!.2f��p�NO�����X	yK��y�K���ݶ�Z��p�s�=���k����QUU%���lο^�e����[n�E�8qŃ�b�{}�gX��	6������l�A�����QZ���+"%5E��2[`Z����R<�dq��� צ�<����38�I�~v(�+[�q���ۊ:ƻ���Ĩ0vj�x^;opX<=Av��� ��w�fwbRJ�����A��]a,���a��M�J�U�g6�@9=��51ib��0�w�}����K����if%c�c�p	�����j���'��������_���a@������_5�l��48�x���+����9�v�t$%&H �5�_$���|�� ��t�xi%���>/�ɥ�(z[�ԉ)�@	[��9��e��_Cy��ٽ���k �}/r)��˚?Nb̠��[�җ������݂�da�5��?$#<<LX!���-eT]�<��4�ʚz|��m�~з�y�9��^8�zd�λ��b�hQ!8�a��`��|/=�X�D�{%��]�ES1wj2SE����el#�V}'J���T3�6a�+d��X��c�E�/˛�*\�m%Ƽ�dG��J�|qEjE�r�d���dF�]�p��ε���PX9�����wV���X89��i������Hى��N�fqb�lFGW�j�e7塚��<�Ϯ<��c�u�J�@g���>���|7?����#!2hgC����R<�X]�(Px��0<���r���F\�I�:y8o�d����g���`���@�����[�NKV#9�E��`�-=�PJ��`j��A%v�:�r<�	� .�W<�8�M\���fŹ1>�Lא�����o�i��&��A��V��e��w�8�#tDE��0�[o���n�[j��x��Mf�iSR���-�NLJ���k��yǩ�>:� uTh �Z4���`Ɗ���<K�y��w�ԩ��D����~��a㲒��v��>3M|P�r�eu e�
�����H*q��Eh������]]������J5���Պ�+gG��Iy#=6 �fD�q?]�U	8F�ێ���]|%YV*&�����h����[���/?����K�&N�uw,�ؿ|IMs�|�����������j��AZM�[[v{fg���{7��o �H�_��,�T(��v����C�!\��\�s�s,a0�w��3x�3�Yj�(R~�C��/������"|H;[��7����gz�� 3;X�_��܇c#?i��~�����m�o����H+I�3�B�:m"�v����T+�7�"W��T�Y�(��}��A2��6#5bQ���+�g�صٝ�-mM��]��ܜ�����`���5��&���ge��>����-eM=A��4{�+�D���9{&��Ӷ�4J��:<^���N;~��YAnS�pzݬ��%>�ʀ�NE�t���*��m�C�V���xlN�W��f����֣�)�u=1##�a
A[�N�?q�&�+f�5��A�/��z=Qĸ�o~c���m�OuSN��F�w˺"˟c�U����������[�m�[�Z��
u��m}�0�@�b�k_Y��)5d8y�Փ�w�=/�s��~l�R��dl$��q7�G�����M��/�&D�vI�T���Q��؊�E��	
E��A�۫�X���w2�f��3m����h$P��� H�4��e�+K�.yF�sq�6�i���kv��q5���qa�e�;m�>zW����/3tJ����UM�Uc��s����+�A�fqZ ���tKcZ� 5 |���MF���P���__�%��q��ߎK�r��o��Ʒ�\e�[@�����lS��?�    IEND�B`�PK   F�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   F�X��) oj /   images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngĻg\S��=�2�
��>zSzG�w�BT���	�����N@z��	��^H'z �����|_�{�?~��疳�.k�}�1TS]��������\IQ���z"�k����Hg����\I�O��ߟo?���I�Е���������:�� ����������ks"OOOk[W��N�<�.��(	Z"���d��x�m�{������O��݇D]kg`%��1�hU�O\dq5�Zl��|�M��l?���c�0*M���Z�ZwN��a��j�ߕ��b���������ad�~���ޒL���~0,�Ƈ�/�7d�|��b)���_N�;��3H�xg���c�AA⿏eri:��>GB��},��i;�w���J����S��E��ٮ����G#�%�ܨ�1T�{���''=���']|޹U��]�b�E�џ?*�������W 
�_@�O㩤0͌����g��A)Z,��m��ąO�s��V��I�k9y&�+����u���58����|������U�J�t�ر�����M��/���;T�1yD2���k�K�%�$Uf�U3�W$��B����K��"T?ϗTa�:�
m�p<k$��W�����YeZ��<[
�7.�����5.����/���y�_���L�܃A����d+�̿��!s��!s
�W�B.�@�r;Ku�&bt�����4��E�Y)!S�!��,�c�����aAX�J����e��[5y���F�,����f�i��x�d!H��y7��<�_�Mv�N�Q椽�Ѹ^y��-9f�q�~�q$�W�
^5?�]�?C��5(��`I�VZ��4[7��|���H��[��S�M�_�ߞ�x"+P�
*w�M�n,5�p�?��}���y{�|y��omj��M�z���4ŉu[_��'u��}�f��!f=�J/��do���{�+��鄩A��bKw��|�1e�&V�~��I<G��t�1[ˉ)$���]w�ޝ�.Γ�Y�"pi�s���O��S���ſ�2�Ϳ6��]�F����n4JF�y0lM�C��!�ު�(�AX�o�֮�Ue3#y����ٓ��2<�`�;�C2�Q��J ����N��c�u^��a�&I�^7 BN��pJ�G��i���q��	�j�tǉ�z*�?v�_� 5�[���W/���)��6mwƌ��%-[���8�.��'7r���xћ!'6^�h �����g��NS��%gvu�sώ��.��7'$���J�L��}�S�/�}ٞf��|�kb�W�)��ء杜�>v�zQ{P�uoQ=�����d�ꃀ��b����uM���պ�X*���`g���s���㍋�G�G]��H +K��,�	��RC�T(��3;��Wτf1j��D�!�%4[l�w&�e+�:��zI�^5x�2y�A�9���7N��e����-i�w���[���P�Ն'lE��)$�ɏ���S��0�a�!m�� �`D1�װ(\o�xoz力�׋��D�߁ԫ]tg�g؜!��C���t6j٤��� ���Z�=_���c#�_Q3��}C ��$����mD�$~�-��I����8 ��Y��3( �s���6q�\�1m�Rc�B���Wu4~��Ū��h��2��z�(|+�q���9�h޷�+9[]�TS�vW��e�Jr@rB�g���/[a�W�1Z��������DeL���O�OyD��u�ԁ%2�(�����{�F��lk��L6M]��8�z��T�B3�x����Ⴑ���gs׉ߙ-�^�6/�r�O�CV�3Z)�]s�P�!:�۟����C��9j��Pa�2��l��j�b���Ml�	��'9E�v7>�o��V�1���u*!�h��ίޕ��	2_G����v����X����D^��l�I�YH����z�����Yr�I����g�}Ӫ�a ��c�Nb�wO�ݝ?j<������Ĵ�ZN�]`�
(��3�i%_�F�s�� H�U\�fz��kw6��w���fË��9}��X�Rx��e�y�d'-�� ��!��;��JL}+�����S�{9<���a�0%��i��U%/�X%��T#��'���䡚��3V�[��)\f�3�H�y�Y<�c��j%��o���vR��F�4�=��K����,�ұ��؃��`�Dim�i��b��nNT�d|@yLV&T�-<��|�K�1��#�����;�W�s�^���]p�髀K�ـO��.���?��� C����kLLH�#N�g��oE��NF���|�e�����!����	�W1E�!G�%�^=;Z�f-2f
�36��.{6N�}�S�;��V�#�A��އ�E7Hx�"t�t�m?<_՟�?��D2AkMb����P�Odv�.r���c�"�x/��|m��A���f�8qr*�����b�u�����W3%^L��[8�Y!Z³kG�7k~ز
�:�S�)
�����l�c\A}�����L�׵�o�Ε��`,���|/��K�G]צ��h�����g���s�f,��4��e2r��Z~�>�Do��6�C|v�g�u뛳��tb�CeOw��]�c���/i�t�L�N��{�7+?�pя�Y�o �W�g���u����&
F�fLd��o^����>�_>�����Ċ�/��Y9dg41���w���:J�B�s��XG��+`�<�vp� �Ê��2�&����!,��nw�P���ك�-�|���n3�{�����w��|:�n�Ȟ��i�~ʑ���;�l�}6)R۹=z��EH4�_��W��'�5���.��A컬�l��_�p�}�����'����ض�Lz�VΥ�/����ƌ���+��J`�hZN¥'ŐS�f�M�ӱMz]Ig�Y�8f��]9M�Ư`�SR�`l���pA����\����u���M��#g�!H���Sy��fm������CO�-�����y��U�&��+@e�Ǐ"R�1�4��T{{����LZ��Z�ж/��}���#U���m����:՞��g��ɫT��k&N�詝O�#z��"{!�زw2�n�r��<8�c�]jǼU6�r��r�>�J@n�W*�U,��|�i	a����˼��oB��~|I�X6�h*k:���݆�Q�G�M��P4d�3s[p�Uk���qc���X��ں���cCs�J�x�-R��tojg:wt��f|�9=�c�a��s��J~�RWs���E{"U�G�����t��tj�*��
��1ũ)��1M���ԫ.=��T�㙫�
����q���H�-u�H�0=¹@ؿW�Y1��JK�:�"��J�\=LJ*',=�g�G_{���I�~l�b��w��G�\��Vk��=�juڡq~�˪��:w�q.��&*XUz�"�Ķ����ι~}kI
�w�2�^��>5u��?5}��%N�*�@R��}1x ���4C+�c�����i�Խ��*/��3����O/܆�7�[_��W�).~b���������72�}_0������-Zluq(���*�Cb(!���G��.8[�~��ɑ'�y�#�N)Sh0��wЦ>��� 9�` 4%�	�m8+������� ��W(��Mlg��f�z��D*�-�ӗ������>t�5t�IO�]�v_w��DA74K��u���^m�1��q�6��xp�'q=%����AP^ݘ�ݸ�nt�t���t7e�Y����^r�]n�b�f��[�¡9�o
����8^հć#n�w4��*�}n(���r���Q��U���i�����8}k㟜o�ש�>y��,�;Ѧ��b�y��]z)�����Zo��n[g4�zٚ��ܖ��i.��[8��L��1�r
&p��{��2���/���k��G�I��%0R�ۘ]� f
�}jY����9�a%�2��]�0�Q�������k|�L��&�Txlʹ>��t�&[Y�ar�}˰�����F��q���L&������;���/WdГ��Z&��N��|�d(j��-b�r�^Cֳ����ܖq��V���|҉u�:>Hf*��e��벤�YZ�3BS�����|JQ��!�6;^G�#�g	>�v����L��yºL_�,N&"�����u�Q����V@�w! �������m�*1�S*,N1�g36�B��J�=2�o����/�
��L��}H�����\��+���������"NwC���-@*�+a���&�({� �����x\!���ԖJfc�ݧ"lL�J�R4ob�.��}���I�d���d{�DB\�l[A.�k�@����0� u�D�	��y�	��	w��[��^'�r���	�ƎިC���Y��B������/���P|��t��y�d��Y���)^6�{�:v@��t$��|�-�&.r��>� �L�zGjv}�	���OgFq��?6jF���)�
��::ߝ�^*���Fz��nOn^�8��W.ǭԂ��0L�:Q�7�<�~���7���t���эh�I��?�@E�?�o���v(:�����5���󼳈UW��P��Ʃ�8��~��h��YN�r�Mi��BNW\D�m}�θ��a�c���������}�)z�l�j���-��1S�;ǣ���л-�`"���$�.�x)xi׵!�rf�:ޗ�vhVLdc2# ������qiݵn��C����7"s�#�Y������lR�+�0)�Cݷj�yK��I���TgҮ�䮇'�a�׭=Z��ўL;⸕*�����@�ƛ�~���-�-&JL�ĺ1�bC�D�r�0�%��~�g\�3���=0�o���=}JEE�ǃ�3����'�/�p""mO�6K��((;;���ar�瓼�B�r���^k�����7���?�\&FIg	|�958*��Jζ̩�GV��!��8�v7�i�P��jɯ��z��p��7}/E�A�W�y����ѭ��D8e�S���1�]t�|v��w�v.`/�Un��;�U�P����2�d�����;tH\R�4l-=l��dZ��(��{��^�-��2��(���0��0��CF���������J�--���޷�_h�M��I�ޭ���y\ ��p�*a�;z�K�G���?S�B@&r��RC˟���v�Z�$�\v^��I�܈n�;[��W'n�~�@7�> �b��4�Kdq��[�2|t����蹃^��6�JRp��@XES#���?G��:�{�*/le�W����yI�u�	�~���VXכ��
����~Үk���['���1_3kO(h��4�Wۍ�$�ac�|�>e�  Ks�����'�c�6w$_p�1���c(�����~Y�u~��i)lG��k��&w��',���B#�ё������m�u��D�!)�]� �>�Z�2�>�fM��-���d+���v�����+��(��S6�X�B����"zLycC�рLm����7�U��0_��l���~hH3��N��JD��1aP���}[z�W�^x�Rt�;��<g��2kS�V�g���W�yꞶ4v�;�\'��w?e�۱�]C��{S���17�Q�L�����	�Ļ�y��\I�y7F�)�uk����X�D7׀K��
�yQ
��ρ��rXpm[[����$|<{�ߟ��:�S- ������� Pe�'|�uF�*:�"�6��h��6��w����:��=1m�ß����-��"7AՕ���Q��/��s���ve+�/JԣM`|��f'��@����� -��͎̀����!�w���'�$�>@:= ����F�Syy�3��D�\	���C�ʒ3�� ?_�U#���g]�L�2��n�~+}��ח8_�o��a*�X5nSD�w��s���g�"��~�i��ްO�mLs���l��}�WyV=�^���(�*��c�Yy� g��'l�Cl�M��X>�U�.�\C��+B���hi	��v����{:&&�[ȭ8UsC�@�L)�P�6VV�<��Bm��y��JߑXXі�`x^Ͳ�Ӑ�~���x5Ke�޳;�F�	"��k�BGJ�,�\� ]���b.�aC�ً.��s�0��r{_��8[� P\ķ���������ʠ��+���f��k�a�ݦ��!Q�⏐
�pAMދr��k�&��%3J�7~�%��f�n���ښ��.HI�U�@`3�[���޷~���9Z������{=��۾�i�9�s����k=<�7���8����;�!�~����\g �D�筕����~^ѧ��{��"�H)l��h��O4~|�n��?��d��a��HU]�A���L�k[�]���_g5&�V�q_�|��S>g뭿��a����U�����9
���vp={��O7���u�ѯrarّ��ѓ��2[%Zmk��_O�l6-2YTD�f�W����g�+�q�w5�~8���8�nD]�V�Gv�3"9�,�M1ar}��m��E����"�{Y���Q����6�U��U�,ܒ�#���t\�dU7�`f��ҫŴ����0Om�e�:77��OC����$W��=����x��{ �X[~�2�f%�8xO�X�[��-ADV9o��D��%#�G�\�3�LR\V�c�N��}������Ís�RuY�\;2Tb�ǚ)��3��V���I��
Q��'���5���F�&
��$'8�f���A��ɄD�ۑs�I'��𻛺ƵVJ�M�?��U��Ǜ'�1Hp�<�Rݠ�U=b_d���)�Rf_�L%|�`�=�]���,�+��G��&��F;5�,�Z�I_X+q�Ln��ޙ�~�|����vT�5�S���v:�P@皂�V�>ݞI,Iٔ�"��%塡ɬXNgh5�w:]ۢ��A��*�*����Z@����H�L�;Jt� ;[ ��4m���N��6y�U���kq���7��������8��3�m?l��'ޞ���j4���g���b��s�U���97�|���`�{���2�1��]L���)�6��k,��Ї�:å�ۂ�<U\*�55F@�3Y�_\T�g DD�a���ɋ�����\^N�.	���^0�^�R�����L�c��9��S��I��}R��ӭ����iX+���~�n��˵�
�/c5pgS�r���9���e2��!�=�#��W��j������r�]|��>Y7�\V����ɪ����[��m�J����u� �r��@�1�6�1�ĦX�<��`�e,2!~d���ex�b��`�ܨu.�{�h	�2�9NN?�'�S^B���wGa���3�9��ɺ��PBo�9�ae�Z�^8�(�``��e� m央�Q�G�T�a��� ܌���Gg]0���^!���k�+�U>�kvWx���l)��&�X>��j��7��e&�<aw L������>��!���S��B�m��G��>!]��ʟ�j�o/�PQxQC
e�/`jS	?;l,07P�5��a�ѽ4���o��#P��bwȂ?[�l�q7P��'H��G@���_nشS�FR�ZJ�[v�vO��q:@��u4��8�3�4�z�f�����\[S��\YCW���0T4z�-�U��J.G�m`
m<����e~LoN4 1�����5��j�pj��#j��x9w�C#SA�����
K-�xN�.�K�i4�o��(��D��٣���K �dP��Ј��{6��@���lʞË�7K��*����@������'������:�*�mp��^���L���Td���
�u� �n{�f�j��)�;�d�4��Ƚ��6MQ4�
AO �|��\ݸ����lD��ig���o���Tk�&�S�q�ǌa_�p��Õ�\����d��aR$�buچ��]q	,ݏ��4�6�5އ555��&`�@��8>�.� ��>�N鮸i���Y2�iP����c��<���p�l��;��&Ӗ��=�	�EB�C+no��Y�ۓ�<����J���*�l��_P�P$j2&Vr62C�ѱ�m�Ĵ�d�ׯmn�~��Ͼd�Y��I�w���H����ۃ�z	ey
�xYH�5AIM�<\�J�Bi�9����SO2���J���u(���U�fC����4�]V�o��������J\xL��j���o��wg���G���tL%A�X
 ��f�-�]E%wa��lq��9�ҿ[���c�]�� 8���I(5��b}c�4����/;8덧�G�џj �~+�6��?�ߜ�,]8�Ձ������U�MTd��;F �$v/?��&t�z\�2@`q�|�?�g�.����Ϸ�Y���j&�%����yԣ�j����F�Zw��C�������c�-[
+�B�aUE�S�<~j!m¦�Wb���j�уy�K�vΎQB�_2���H�`�|mh�:�^���zA�Զ���f��Q4������|���<Wj�o#���zNm&��	ͭۻ�k�����o�x�=��N�pz:9�9Jh5�=����&H��z\�����X��1��������s�S�rkF�	K4?��c����]ߜ��˝��v\���ޙ7s�\���#
I��SSu/�7V37�f��ǣ	���	�U,|'Y��8kd?W����������+ ��6"�]o:<�]�6E���+류�I�q@h���Y���{(U-�ʤ�ؗ�.��R�C��q�s�e���"�xr��/�<X��.VΞ�6�����|����%�\
Ҿ	� ��O�����Te�X��9��%��x��녔n�i[�)���El��4�����[��u��ae
�SVSX9��<�Ǉ��,��	{n48$��K�T�G.�D{{�k�����k�mG;��F��|��2i�m��r!��N��2����.��?-�a�C�s�,�d9��y���G�r��6ڼ�>:w�:�	`��H�Y����l��#��zxdZn�Ď�y��X�:/��&���%��0��<X����RW����s�yK���L[Q��/�ϛ4�6�-_�4W��蓡B�>�ΰ��۬��O�QI7v��fKh$�be�����ٺp��z�����WA�)�����vH�h'������2�bz8�F�Y\
���wv�j+ʗ��LM��K�<d��l	�j��ى��C���&�W52�"�J"B�'�*-(��tR�����р�L���5�"�~�'UjZ��j1|9o��dT�T� F���P��`���.��e^O��Lk���w^;�>�*�=�b�����+Qn�N����Z����&#_��oV/��۩���νKZWrB�A ���w�b��I8{=I2�Bh�MM+��vu���8A�ˉ{�δƓ��!I��풴| e��U�{��Z�£+��@��o��B< ���H���K�s+��R/pn�@�-��cִ��\W:�W�x����=��e�1�g��Y1~���e�$'=~����L|�d�|�~�/����/��̘V[�kmCKe���r}s��_ӥi���+�م�Z2H����v�ϒf���g���b�V��0���H���ݠ�H`R�`9���ۏM�o�z���,U��%G\Jt[�:�Ӧѣ�e5�0�{�Oj����7OJw�u��8}D�X��(?�d&���{���`.ğ>�;��Q}�f3ͣ���&.)��#����+5.�J�A=�o��o&��,V���Uߘ��5*5i�`%��v��z�;Y���C�Nf�D��{�SV9w.u�������ĝ�����f>B���^��c�����!�n���O�*��%8�UO�������S�'��6H�,uO��rG��.]�t*����a�_8����ky��j�琎�
��7�\���/����_*� �o\ҥϊ�s���xr���!U���0��������,�`�.(���A8��H��B��*<����]2v���f�R���t����*�
wqO�F\H_��I��R�;W&�g�	Cq�,|���U&�f�=�"�݁��W13(�����=����!*�z�h�I����Cac�Ϋ�m�C��3	�Y{��@]���u���������LWZ���p��Yc��;��|@l����*�/�*VC�v��[��)Z�`�ӝ]��y���׏�ofl��e5��d)����PJ2���󰜙0���Y�Mݳ0��YQ���㟀�^b���|j888X�ZJ��&s���x�P��b!f&w��a�`��	v���}��](�q��<Sx��t�-��
��*�QU˲�]��ˊ����W@��dq�]ۇ�������N��T��ap����4a{$#��ʵ��#�XP�<$���#\@�8�-o=eT
���Ĳ�C��FNx+�+֓}�)&�M��/���8�ш+�X�����!$j�=��{�G^�_ NN�~{5���R| Zvg��	��Q�3�h.X=Lf���ߌ����lQ�=��O��ٚ�/o=���ӳY��,	�g���s���3�M;S3�*�9bS�i�>�OH����3S�Q��R%�vdw�1PX�.����oD�D���a�,�g��l��U��IF����5 ��}N�!�R�V��Չ%��c�$Se���Xy��i�}B颋m.��� d�2U�m���#�)s%�}���ˏ�O=�u~�z����=�81�$�1F�P̳267�3Se��1�,����0��'����䖅����D|�(�l�?�f6�1�����>(p�.����1E$G�<A���p$���t�����w���QNr�nAY��s�I�Q�)A���������F��i��q�H�\+�wi%9n�'qU��%_:�d鍋;W�c�?�q�5Y����k���c	۷����t5ޜ�s ����H��bH���Ÿ�.���Ƈ2�x=��zV$!�{C�r�y�� \��<��{c�_dT���	°�ժ;�py��顺��.)��םO��b̊�V�Yn�Z��0Wre#b$N�k6-�+3��?��%�*��d�!8UH]�w���z�ґ�Q�L�a��$�T�A}����E�\ �Xx����?C؁����bM@:�}����͚<�/����`d,W��(��^:�s�	i�V7�1e�\�c�l��G�
�˰𓾰&��{Ҁ�q����^�48}:���j�=���X���3�ڴ޳����:l[���w�o-]�����i�-T7f�{�t��~�M@g�L���ä������+���(�u�fվ��2[^օ���{d�Y"�0����I����!(��P���|�IҠ	���R���o�~�Q��,�4~a�c5
R$�;�{������Mռ�u�����Z5G�xE�������a�/�?W�UIy�#����@]Vb�����B�OK� �/�����6�ɺ��<x�d�@ �Q��k
�Nv.��6�Ȇ�r��t�۽؆��u�*6�YU�_fk��������C����Q+����6�ɾH��6=��Ǿ���'3rvWk��x��O�.���{,��{�G%��C{.���VF����{� :��_ʨ�J�#oPo0���[��HY\��i|(d��+��8��D'�PKk�Gٍ�jl0����2�ڱ���a�C��Z�km���&�}Z�?��v2�>���߼
~��5��g�;�#P��M	+�1���9��z$?"����΃�M��/��4�{�*.�Ѐ�����>�S���W��I�wy�r���y�^�M�K2 �NP�q��!�Th��͟X);��ʗ�H�`�<ᐾ�[�i��'f^�#�R}z�(���/kE��)7��$��ׅ<��[)�
�֍CJ֖��'��5�3�j�lPs��K��V��aO���l��YO�|��O|r�5Ua; �H�-z�a&�W�sH1�	+�#&~A)�m+�vD�%�U}��z�mN�u)�z}�l��
K=o��_�_�?�OX|��ǋ�`��ir��$�c�]���_����k#��h'���	�eS�e���nB���4�&#1Vۍ˶��I��p��ں4GIC�kc���C��c��8'��b���`k���������F���.!��N�vM�r��v�\>�Ą�7��M���w�Y�f��v}��Sb�'V���͒xp�!�2xUU����a�~V����gxX�.5�S�?����r�5~)��֪%�]{�+鼘�7Ӽ?�Z����G)iTOb������������(.Y��ŋ���P��dڬ�n��{-�	cݜ3��Z��3�:r��S��G��2#W��
��jk9nF�Qc9��lR�]�����[{Ψ�z�?���]4|p2��`EMbI5�B�+7u��fɝWР&'iֳ�7���bl�����<L�E\#h^=��B�����_��;���^Y�)`��6d����֕^����r-*�j�)��p����ϔfH}=uH-����2Ϲ�$&�Y�x}��\j�F�c?ơw�qP��nq��/���P�fs]��.����ݞ�q῁Qӿ�;'�&t���o��y���6���|��X�p�1C�އ�K���9mK�����P=���}_/�� �u(�8/ƼmNV���t�D��d�ed2M�k�0���O�N�)�ք� �ɫ�k���Q���M���js	�vU��7��b��4Ԟ���#
�Gt�B]��o�0OOx���M{_�3tw_��w�`�>v��/w�it���J�N?�2���	�Zi|�:FR�����7`Z`��?���*�Zn��F��~a����{8�X����=]��#zh>�����Ԋ���b�Yj�#�����g
.�RQkB?.����|���]p�g<�����֓�׬_	T������2b!C�E���x	�^�U��/���m�j22gՕE�����]�B?�B%��J�$�j�����,�`���}�4����<ӎ�Z���&O�k*TՈI�] ��Ӟֵ�/XA�=�[�`VN��f�"<���S���ه��b�w��`2��.�X�7�Rm�V͑�Qn����V��x�G�������o����z���|��I�?�(�ܙ��¯t��OΟ/h�ǻmZ�.���j���?���*�%�ʟ�4L�.#���RVE�s)77Y�s9����? �io���X��%�-���x;q�p�ˣA�ҋ��v)?
)᧻����Z6V0��\��;k�( �x* ;NvT��_?=��^3�xЋ�*
 (��(��m0��V�1���)�G�;�Տ<���t��'�m�����a]�|�hq^�N�	8%���Q��Ur�SF�=J1�p���H�0��m���o[5sg[�0������_���^�뽿�_RV��u��	?D��U\���_i���N�0�v3�o� ��~�ɼ�
AR�;�]�n��?���
S�N�\�
�vt.P���+K��?�_�xnb��,ȹ���b�;y��f�����Uǀ7��.���(����HQ����ôh#>b��u]L��a�/��fx��"��L��<��i�!N�e���X��2>� ��V:��3v��QB<���������A��z����!!o�X�\��_hPIE��Ѐ0��}��Gf^}��%��~�W}D�v��t����#vy�Rh�?_e�*�Uv�8Πƞⵝ&1S�6��D���n�$��F2�׳�Gقz:q9��k�3�:�}9Φ��>fmL�M@�V8̏_*U���?�;�nK^��y�-֤�-�:	h>,�w�K�Z ���}iwǡ4Q
u�K���%�"j&��t��O
�6�����v=�8���]\S�HŔ��[xzڂ��[ג�H�$?�Hz+��$����÷�}yt���WC����ؾf�^E�+��Ÿ�j��d���i�]�I/j:>�H�����3�B�a?���ۇ/z�k�:M����N}'���6�<�M{�H���x���.;B/�r"��l������O�c�/�H5OqzJ;�|�bSN��#��0ʺ����z}3�6Y��y���\��:�L�Ld�O__j\W����"WWwwrt�"��3�B�����_V���bV�Rb�Ѽ����)����az,[]`���s�}��$>~E�R�=��=3�޴���/~V��e�g�F>��]��'�MM���Y�|����^ѧ�Yeoʸ:iA}l�OO���~�uB�9_�ڊ
�r����I����ݐ�<��'�w�n��?���=�}�U���EH�%^�D�4-L��NS�%�Dg�T~��6���b��rl�ê1]����R�5/G�#�O���B��vy/��K���ϓ�|+���S65m�!�37�S���S�,�3z�
4p�Q�]��!�o���1��-n�IW)�g��'�|���'������{<��W�U'���K�1���k���kc By���� ���KW��ge[ճW����=�WQ�e�M����Ǽ'�Q��S�����mUe���@�+��ѭл俆�㲲�߸qC�g�q�h��o�ݏ�%��Q}.�T{�
�6�R��|�yk#1#����c�W����.f���Qr~�����}w;�n��\$���=�*��`�2���C�-��x�:)OjiTd�"�>,�}�_H�����p��|�������~V8o�6�^�u��ߵ9�~�
m�=�Xn�Pm��q2xp��h�霺�t�-��}_�}<;"�W��$�bl�q��-�E�dcs�rb`\�󮔺����8���^B�f�.�Ul�,�>�����{���\�ԛ���U�%=Î�`w�zGH��=����8\�2�?cgz�Nã�tx���_i(��ݩ��g�S�� �τ�+�;���P�	n]�ҧ_��6N�9a)!�mu���k��{ɾQK���ڗȑ��DP���#��I�^��b���T�{�Q��[ʥΟK�d��	�h�?���5T{,L	�N�GG~�brS�\��w�xyҼ�_�����F�u��4~�	W�A>�����R)�_ZM|Y���x��D��4��C���N�>�S�ӛ���.���wo'�<[��|֥]��ǁ���<M=�[)�ܙ��.4`L|�N���U��-�Z�Bҹ:{�TGa|�e��������vά�])�:]r�p��3.3�3u=>� ��{_,0����&fͻ˞��&%�/�����!��������D��o��a���)���q���j4����	���l�u�$fZ�_�+���eRW�|�������0�����sc	��Gb&g�q��3�t�򛿼�Wi�7�E�b��$��;���r�U�b��{�*Skrپ\�m��i�u�.'>�0�b	����',>�0�E6�|W���6�P��#�[�%4�O����yX�����2>k�D�<�����uўs�
?�.��-�����t>x�h��rҴ��a�f�)HY�o���;�
ϑx"U�^Ys�H�;�-����C�<Ðk�B\VKF�Ya�]j�u��t+��H1|��i�<v$�]4��S��U�P�9WH�?sn������5�_����bO��~�n�r��jF?�_p�`ۈ0i,w���`[%�����������r�vڤ��y7F.�Ky�N?��c;�^��D����<�� �k�t��}gZ|
���vv�8����߅"���N�_�^��b4j.42��c7h��CL5��K;�ɣ8�w?�u;btK}*��O)\цBu�c��cz�o*N\�ku�������3��F4�?)���ԇM�f�D��O润��')>ʴ�x{5���뫍W�4��nL?�tq��#�6�i�xy���49�}pP��^�+f?]#u\���s��a�1R��'����x�~ay",�e��g̶�'���;[�S��{Mo�ɀ�df'���C�\ӆ}J7�����Ơ){��[߲l)4�s��'��)��UA��ύ@��JAb
����b�
2�ѓ����q�:oi^��y%���q�V���3�Xv�n�^��_��-�1�!���͸��^�P���e��V����n)(�r��w�k]|t�mdP��>/X74B[;ܾ���	@� z�z.Df�}݁Q���n��IA�Lg;�����0܀�9�w�W�X��%#jv������C�aS\�f�������hi(ɯ�Q�5��6$)4�|~��su}r����Z���<r������י-g��F��_B;v20�ߚlK��E
>.�wS��?}�,� :0Z�}4�� �\��)>�o������q�㤥U���<�fX��¨�K��[r��S꘥�ƶ+-��1:�s}����h�(>����1��P'��wa�s�����q-�JӍ��uy�t8���$HX��x�P�o�7�k�U*��t)5�o=�#���Uǘ{������^dOB`n�����3\�� �ڶ�uZ�v������9���c���w��Mn�
�J͸����]܆
��^��7��L���]�f���n���C�[��
���!K�����C�y�|]|�������ѩ�z�5�.�ů5]̆w�)��[�xa��&i�[=����vW��[�ǔ)�{�LX�������\��M{�_�=�sx����F����5��!��]�ݤ�>S~�K^��u3r69��5ɫ6�E=����mv�[r��V+#1_#7�����J�1�,�UFD�ȳ8�ͨgs���=&&�}|�9�w;�Ь�ƽ�A��hR�K-�n���E����,���Em��e͘O�>P����{�Ze��?���q�<���(���f�q0�KV��Q2�����]1'3��K24������$�*6�c"V��\�SέkG�-wwhQӒ�����xX4�,��V���Ӎ��Am^��D���_yVj����}��O[,��1%�@q��Ɩ�Aa��Q_�����y�;~�_,
/�(8�|@`7L��PW��@��;&w��^t#���,��<(��h(G?4y
�7����Lb�I��S�7��(�_+Z���F�0\�ch���z�xc�=���k�$���k�����&�A�CB���A������S	��;�����Y�ߢ���;���0�����\׉*�ݒ��ް⛹6gv���5D�bO�!OҜB�߯�ԐT�B�\߽�l�ȢW�[�Q8���Zk].�p� ���\"�G|Q>~��s���C���Ć.�tD��;����.t����\|������d%N2��4����WxG��]�7B�_���4~���ax���!��BZF�}U#����wϊ7ڊ��s��wM��[NԵ(ԤiT_��4�$���Cr;����b�W�������B���?m�/�{��'Pܕ6��~e�H��{�۟_��L�Gpۂ�Z[��z�YD µz�hT㲷]���b�v�Ma�T�M�9���C��C�@��c��J�KY��yH��x��-�h�\����˒��m�8�r&����~�ގ�j�G�*�d�qB��'^޺�M�X�y�f�Jg���-y�l��5��_���UxU��9M<�	�f��c�4���I�V�!V����`��"�B>ka�-������%LȬ�h�S`b51ӥ�y�7;�FZ\�
�#.�S��Q2�� Y�k�>���@�E�����__���}.���Z��{+�:��
!W���͙�(�r�Z�0�^J�����/\[P��h�lR?M�
ZB䑬9��8Y�ۚ��w}��E>�3����x�8�81��wQnn�i䷱u�����z޵�3�Bp�Z\��e�RP�0�tw���8�y�t���K����7 G����x����)�p��B�q� g�;������������Rg��7�w*�]��!���?��E	_��t���j|R���	��q^�6o��SΘm�5��r�(<M`�o�s�r�!�9&6��N����+�{Ƃ��K��N��Y��5�CfL��Θ�G������b��&��]������qO6��GƧ����e���U�ϕX\��>R���p�NW$M��T������>���ړ��L��@؅�d$���Δ�Ҥ:W\Y�4��m�v�|`�[�l�is��)��*�^�����+x���%<%g��{����D	v����Y��5!���Vk|>��c�?�q�J�I�q쩕�㶉%���������^�*a5h֨}u��)k�yc����0kv������ <�$-8�~��پ�9ލ@or�8�fCH*�l�]������`���1+L�xk��M��u�o����.����?���8��w��m��*.�k��	��[*�*R�������v���bv�Lm\�v�	��熥����wϖ�ֽ�gZ-�M&x��*�̹�9m�e�.Q��$��l4�Up<v�f�4ġ�"_F���-�)v֑2�C���/,��0�������zRy�ɩh�6'\5�U�V����IV��!��@�����l����Y$+��`�ݪ���{�(M��Ϙw�wk��ri
��~��K�����\���T�����v�cf����e`��D�\�5�I��z�������8�{�co,E]�<��o����S�X��]_%�_���$����D��f���̂�L�` ��?��з�����S\�d��n���ߛ� Y����*6h@/�{m�-!J��~�
5l����g�m��ւ�c�7��[|&���ה�isC^I���f���}�#�hHVr�1w��zgf�(Y����5uUf����K���q�K����u7n"�V��}y�y�}!�'��������4��p-wخq7ܬ�S��&އ]�UP�~
I���x�jC3�z'��y"9&�Lb��e�V]�]�

���$(l]Pm�ē*t����sw�ur���(+W���M��*|.KMQL�@H�ztw7R��j���mӹ��Uƹ+�K�|t
@��t ;��,'� �n��2ŬKZ�kL�=��th�L��\嶕tt������%[�������VnR,�'�q�)�̟���u(���b�/�����sr�U_K�(��~3*1�z�v��l��c�s����o�|6)�~a<�Z�F¤������0����Q��3����鷙ߪ�1�(���A~��B>�"�~2�[.onU���;~\ƭ���u�Ga��l)d8��ψ�I�Pۖt���\�3;����r���vb8m�7*����Bzi�>�4�Ĺ	�65����hZ�AZ�ڑ�#����ר��n�KJQ���/ú�1O�'F���!������ �781,��.y���F��:S�"(����8>�����''��-��3��Jv"	�k�ר�֗6�.Y�7�>/E�N�Cg�&��9)M�h����L��[e5���q����?�F! �<�g��c⡸c;>Nd|�:R��x��"�+Y
�	kƬ!�����k��n�޵����-�?�;�@�ԭ��k3�x�ѻ>��u����b"Ԩ?��q�3H:rݷ�upq��È�����x���u�`{��`���q�:���he��+�Ն�,u��c5�,��US*�Ō�=�r�0��L���љ�N�֮��/�o�"����� ^f�]�q�-f�tl���5�� CM��M�NET�Q��T|#c���@FN�|4�O7��QDDDp��gL���=��gޛ�I�ȵ"7a������%aI��2��O6���gغ����a;�U�9���Q̏If̋��|���n#�}�Fϰ�%W]��m,U\���׿�������mV@O[��é���g�����D��D�wEBӿ�/�`��A�G������K8PgS�(�}��)��..�Ws�^������[��s*��q.[�����	����ݮ�b�cB��Ҋ	�>6����]ە$���N�[�Ǽqm4�#0�S��Y�ed�44�rhY���*�"2;���	�Ф������Cea�}�aRO��a�0�F��:X?�s��R�?i^�9�����@
,{$�z������S��rDiހ(�D���50w����N%�hE2@g��2Эwa�!�n�wΟ/	eu�ܹ��_��O�+�cBvU���/��1ש�_�;�� ��<d���/����g�V���Xr���&���У�������M	�6D���.��ll0��C{�?竭b҅���G��-7:�4�?u����S�ɷ����HQ� ʄx�|Z&u$EY�TN}ϰ�CRB��]̬�ٵ|�&lw�vK�S�6�k�zʁ�r��1vG��eҘ!T��ӑ�ɞ3����Q=��!B�nZ��vZ~bL�ro�q�v]]]$����3���M^%��{X��v�������)���k���}/��z�G�Z�4fu�p���72�]��/ ��'�Xu#3�P�)/q7�6�"k*E5��/p���Gb���9�y'~IE}���:X���ڨ����;��X�W��f�p�ՙ{~rZIӷU�j��)�J51�;mo\o��R2�Y�{�xR�V�����d�YWiQ��vZ���F�]頃�UB)��ue�m���!ϚC!X9Z��3c�y�?;�r��;4���o�gN��ܔ2�T��?63���-uBu�����*��mG�����r���
��e6��)ϑٴ����ǂ�F����|���]8��%`K�%��ђ[�O�V���^'���8���w �J��Ȧ��3*��@�S������RD���� �˒6+u�����T@�%2�YC4\M��񢢖IJ��C��\��e5a��,q��]�{f������&=�����*\�/�1y������Nx�sVjZ�:2a"����A��ba���|����� � ��UQYp����r�������S���[�.2b1��;e�M��{q��z=ߟ�a�l��*��^^���׶Kx9Ԉ���W����$�������������KҶ���M+�����.��p:�&\o��e�?�����|1�?���A�|��(�ZP[��P#hځ�c_���ٌ���ռ��a+���ֲ�?��!<ɋU����D����Ђ��p˛����kt�a�ㆵʤ��R�,��H�	��Z��8����g)�)���JOx�P���n1��ف&�$)Vof6��+�A܎�?��|�P�2���ԋ+�n�Kˊ�^��/�_�j�}�S!'P!�Xϟp)�tw�Q��Cx�S�d�j$��i���㝺�h��N��� �Y������ۏ�m,�a.=��N<�XЌ0�54�}����{�L6�І�Q�^_M�\Z׿$|��;}��N�0C��,^͋�k�C zgW���5�)�j���fl-$Z3y�(tFT��k���!�h�2&{�9-2�����1'C�CE��u�|��gE��x2	"�J)���u��Ξ��;C�Y��{'|l={�,�������%7�Q�c#˽F�9cw���kɅR��/��!Rsoǹ�/�&ٳ��!\��X�#��f,z�s���/�Y���6�5u/:�[4�,�����E��-�.��d��e�J[�ߓ��܂^b��O������:y:���O�OgU�#���f���4��"�݂�|�|�7Vi���w.`6!߫�rl�m��賬�{�bI��"sB�y�hȆ$�?�����"(�޼TBA]`�X��/���,b�	=�:iq5���c��hږ I���y^� ��)�}�^���?���L^��zv0�z�DN�<{9vv��Y���u�aP�ƀ���tdѝ�1��ތ5�(\��?�h�C3g�sM�$��C?a���
��|��hG����{߿
���������w�w�fo7�<�U��d=~�r�V6�i�� �V�c�j�^#�#�C�
�ʑeJ2�r&����n���1�'`��z,]��A�a���5ݜs^U-|_�G��b�p��y)��l�4�&�B2�iQ����9}!pS���O��=�Q���Xn�D��,��o�z�[�]TRs>����z��/U�����+ދ�>�������ן�8�ޙIƸPK,�3P�#�1�m�i��=?�H���"�lXC�O��R�x��8�����v�_���<���:<I-��2J��^e�(�O:a��;$8�:�p�:h�+��<o�C:f�,���:W��;a�t]I#���A��{C�/��й\mnY"��0w[: ?�s}�9�,����.J/	����%����ӵ0\��WN״��ǿ�^q�6;D��Y���/�9����>q�R�����y�UJl9[���R�B�L��X�~%o�Pgi�t���;{Є	�O%nud�ʲdn��6iC'�c/��n��g�&^}_������8�/&���(X�����2�H�Ȼ\�O)����y�1y�|���C"��eq�L�5S�������.�����?yx�Qq���h��d�Ui6p]N�mQd��o_1z����+�vYJ�0�u�[�i����6<)���G�2v���� ��`2O�ڃ���bÎW� �F�y��&�t��DP��c��Q~2�rDkb�͞^gy�Г4Ѝ�*���'�[�"�����G�����@=���܌��D��6uT�����z�v��W�>��_�$���IY�_�~�P���>`�u�p\����&�v����%ܶÇw .�|̃9�~�cBw��U6|�,�a��ئXWx�f���(��>݄�gOl�c�wO����ݮ�&QaEY�l�!��k��?[u+O�A����Vv���%C��Y���'���1AA���^$%{�W`���sR� 6���hpm���H�m:����j�-�j��?���dz�;�#��|�j��ZAp�!�FB���z��3�
�
ae��fUb�z9�b������S�cd!ۛ`���<�v��=��g�#�.�n�f[�OΙ7u�G�f�.��#x��=��������&�*�+ⴠa�opa�,Kp�E��m��ߴr<��8r r�SY�\��tn�����7��v�@���~�_�4�����֊<���3̒��WPN��'1c4
1��TҎP�Vf�]��o�'-;�gw�p�с��|��_�nY�}0~hRme����ѴHڢ�4� �ǭ0~{H��/�|1a�X/��(��T�I�s � �
1?�k=04i@����]~ƚ�n�,y۾/t�V�f6�.<��_a������-�z2��5���SI�Zx�z���L%�0Zx��%��F<���;��9���� ĩq��J=P:K�$�|V�b��z�6v}%�ni���X '�~Bp�.��'{��e.ᡝ��{|���e��e)3�x��SY����HWb�u^*��|mJ/��ǣ빅�53T��cc"�Y�RQ�!�0��t�!�-��<b�"�]0��_.�9��^�֯'��$c�^�u$��)l?�IN�5�?��.M�S-��ȣ7��Y�H(��9�01���M��:	�c�����%��Ҙ�h������a=� �[��߽l}%f�(kF�q��P�hq��f{. �M��d��"|- �/�k���-Ccq����(h���W�A����`(Pvu-B�a�k�Hxۻx 	_��+<2B��ٿХ���"G,������>��n�k�ׄ�*�ί�0���U�0�dwz�BH�?�-j#��rr���/�C���}�&{�㵡c;hB�	��tȣ���0a���\f�L�܎�Ƈf�A:�=;=3�������>�4�9�.fgl"�f�x��賛o�ۙ�F�~��-J��F�>�6	���T�����B�4n<$�_=+YF��\GxN�L����pUPЁ����p�����>~�8|�j�,L���~�^aS4YƆ�����'�֡�Dg��3�WHX�^����Y3�[n��1�"n#+�Z��׎��H�(��d�dYfb��2	��&��u���Ls�i��1)Vzd�2�s��d��/�>͸ل���r�0��z�������������F�9�5P�~ʟ%&��{р�{�Ӣ�˥}��~�4�u�8tI�U$����~�m+�-�� òh�/�<.1)���JT���L�P��|gRAv����m���"�m:x.l�B$b4:��t��x^�K�	q��]>�Z颎�/w�g����̩U)���Ƨ#�U�17R��Loj��/mz��YG�������\/�N.����ӻ۝����K������zOd������￉�%�M}�Q�p�O/�k�����A��u�6o�g����~T�a�N�VI�b��"�Od;�Ϯ� �w�A�G��d�����/��ߠ�F2IA{��V�2�n���jtzU�{8*�2������iK�%J}���{2�{g�#�@u܋�/�'���)s���d-����.����V�д�����ZM�9!<:P��t�>=�w'����A��P�� �D����R���d�k�
��31�ܸ7�"c�/�G��TbĬ*m^�R�}y^��LL��f�'K�И�94�P��"�\��j�O�_�>��a��tbJƄ� ��Ij7�t��@�ko;�pZ٢�6�*56$�����*�U5�|�O�o���5��m\���<��s�5��n�?2�Ni����EG��h}�|�����3�)A�/Q���Ң>���6 �l�tx�1$�}������c��IsL&H�A�"Hj��5�7&��o7J;.��;q���M�2ǧ��{�USB��'�O�)� �L�Љs�ۓ7�I�����d=�.�d�����5�c����ِc��c�7�8�Kē8�\}�����s�ګdA5`���8�c?���>�cxJ�s�6��e"�_�$��ޕ����Q�Z
8u��Z�'-��J�#z{%S*�0����M���ӕ�/�6�4wuf�툦s@)I��/�{�	�)�z2�S�j�^��d��\~��A: ��$ʺ��׹��tX���l ~�]��\�}F� �ǚt��6�;�V�xED��8%��g(�Y�Puul�S�������&8�ݜm�2�0�N�vm"�V,���r�L��u��]�Ѿ�&�\�ox�O���Vj_�|k����$	'E[�$���@<�E� ��8���H6ϕBl==���O ���I+[�LAG���s�=��;��R�	p�f\���_�k4a����bu����M��6}~M<Zo��T *L����ex���gT|<+&�v���-��(��0n���$����W��"%�'1~I��bB�ܑ��/Jb�N/h�ܭ��˿�uzˊ�uS�!0qh�i&f�"N��=��5H��K��6a��B��=����u�I�͐!��X8N�p�ȳy���!ȋ�Ȅ �
)44�&?�c���z����+�7��.�y�c�x�� ��j�����H���5vu�t��0\��\�5�_p�,4U�l�P��t
���(Y�1��{��C�S�Ab�G��5{���͑�1�r���$�'Lں$�b��s�v�a���H{y��/7R3�k���ٸ���>R,a�M�8#un�D�Ӳ)ta�-, 9�:0�����U\ܧ�:��C%���M?�$M\?i����u�˛�{wD܇-���C����giX������v�Mޑ�GC�����2%�W��m�G��XnaGiޚI&�b��2^vE&�P�r�dn�A��":�u�gJ�f���q	���q��.~��fQ���ĲTZ�r��e.Ј�LB�e��Tv�C���7��ں0���|=��s���.�.$E��T��z��vӕ~�����q�=��A��v1E��[�g��\�&�̐6	F�_���Y�Bs4{/"|�x+5��R��*�!B�4�Q��l1aP�s�>@<�����^S�gS˔�TH�cD,�'�ٙ��^��ۿ�r/;�?v%	�a��Ļ��t_�z�^�E�%����+��\��'�
1�JN�R�����Ј���o���yqWG�&� �ԥL��)7[�g���P9�k���'�ع]��6R��H؀:\VD��s�` �[D+�+ށxc_:.^�jAPƅ��$��*h܁,{� Us�W�u�-�V�~�!q����G�N��{�9	h���u�ϕW*��YHrH�m�PU�I2�}���^6��m�9��T/!����o��=�0���bb7C�����j�� u��lO�3\!��M� O3uu\g����d _��O�P
��40���&���9B�P ��w����㦃���R�|{�^Ts�qb�CF�B%z�_h��1R6�O������OH��3g���1]WPx�n�JLsH����Bs��[��/~��X ]�L��<� �0^��vk����[�3��(���R��E��}^VCYi����c����N��I�(���`߬'eX�FB������m�sm��*��ݟ+�Cʃ��uSG����S��q���_�L{�����ڸ�["�ڤg�=½=��~�Ed���J�/i�ArT�_�Z34Dθ��:e��8w,ͬj�AN��p�_.�Q�㊾6q�,s9����}�>�
KOW��v C��*Ѫ�Z1"p�KK����Xz|v�����A(qݒ���T����o" ,����r�;���$$R�T��4� o��IxD�u�2�Um��ԗX+���������fP(S�)�e=�:�P�sqK��K��vO\*���#�k>�(�X X�h�?=|��O���\<��ת8����М��.�D��fV=CS����e[��e�ӡ�	���j���b��y��[�MD2V�^�����yS��-�R�V�oS�jD$���R������q�s��	�ԉ���:0.��b�\�OK�9�Z��ؖ��'�F�R���N4}�RtS�d�.tiGS����~��v�Jf��=s;��!Y/o[�����=�l���n�C7�W#V���U��Rn�l�W�+e���(1���2�ٕw9��"���V�V%1��!ʯԚ�k�A:�%j�g��J3w�@����a�5��ް1�2/�1���g�ʹ�.�KLKl�drKg1�`詸TL�D5�M��᫺��&D�&�m�g���뜀(���L�4QJ:;!���|�F��6k�d���IF閂H �'R�p��;�#ƪD�����6#7Z67��l68�y�\��F��Y[�~W��l�)<�V�9c��3}IL�w��R��� b^"pfs���Ȳ(�j~7��XѠ7OkRydP��F-����g��Z�	��<�K+_��s��av��3'6��X-���c&�ٺ�o����ς���������'��y�\�@h5��Gp.>����lO-W諴~	A.TMWπ9M��Q�yU
�%������N�+S�g�	��$s=FH@~���(+P5���8��|U���?�_*�0n�����8$�����-@��$��@S�����}�e��ˠD;ٴ턄-{�����1��M��GtK �U��%����h�
I�M�u�\d'���3Z*`C�܁T�j�%�&��܇��Yf���;�9.$oE����gR<-�}���b���W �c*(�rE�zH�r7�팍�"y�`��,���%/���I��:zv���r���?$2�6c���h�w��=
���~|'�'P�9<��]�.�O�}7�|}����̄�v"���Y�LO�J��i�����b��lL��۰�NH/�MH�GW�>�{#�G�| �;V��.��BqA��Ͳ.\��B�%9�����*f4�8�8�!3�V���p�ӧ��HHrkI�2������҂�NCۛ_w��xW6�$�3$v�ǩ��֤�bq�%!1ŽWw���Sc��� ��n�G�#veDl�縋��P��2�/ӝ*���EQ���TH *Q���C��
�XL���@QI35)�q��,���,v���C�:����Ͽ��܃��`����8p�+�tsm�f��b֦j�D�&lS��'K��MU�ޅ�rUWk�5m&��4��-9즾�oι�H�Lzh߮�E���K���CPVu�z�JG��F4�a����,q�����'�צX=�d�?�OvCY������8ֳ�6��e�~�n��A�����M���>��v���啊��SHy�Z�̈���C��!�g�KT�<%����(��I1Զ�o����˸!�4D�f�):0�(�b�*��W(C��9��f[5��J1�p�Q��Ыk���JZ��]�g2ޚF=�<���ް��4���Eڈ��'��7{��w�D�O~���x�M[��0�囩`�>�+��"�c>W�2�v�c�k��3�J��Y�� D���Q��  �ާĦ}��\��m6�`Ӽ�V^� �1�D�g�ȳȦ��+<x�(���N���W�gKR,0�d�멏���r�mP����q��.C�z�hX{3Q!R�Ik�-�<��`��Ξ�>W��5ڤ�:��˥+��U:���pħGj&;$�#^���I��^+Nr'�����Bu������o"X[x�h�iu�8̒b�eBu.�^I�k���?[h����J0�o:��h�:D;@�S �k�9�Ci5U^�D�ӻ����R�qɆ����ܽ7��\[��a��E�^<�Rj�.�u7pٌYV���mL?�z���aw�{J%Y��_��;?f�����@˧�+���uF1O����|�g!:-X���2ESr~a����.s1Ze�k�ͬuC�^�&l���+�^���Z�X]�<���D`�X^��ћbw��{�$s��9 M�xAD��~��(���)�QJ����o�
�Ǹ0����>d�E�W8�7M��#��2idq18�)�k��(��x������V: �0 4tC\�
e9R'�{I2X��"��𑠗.���"
1�a%���Lt�/P8���p�w��@N���n(ԍ��5�ڞ0�z���3	�$D�����4���Q��҃��o���w3kC�Ó����6S����jJF/�A�ɞF��=\K�Gn�G�"%�W^Gb���]<�W ���lP��F�zs��bi��e8V~��Jt��y(����p��l�t��+���Ѷ�_�k�IS&O�� �uȦ�I{��2�Nj��LS��+���W�q�\G�J��I��99�6�{�C79��&|����������/Q�9ċԂ�!Z)m�/K�xe�8Q�%��%ҺĹ�!Wx�ʴ�
8��J�=���%���h(K(��2,J�Z������\K��4���_},u/VV��!	�G�ͬ�����8] ��f�e(��P76d�Z' R[PҪ�D�X�J'�KA�\w*���+�\�@�l�\�SϻZ�/�8b;���Y���?�����,��(�R*K�6\�79�m�Glv$i!�����5�bȿ�(��GKD�{�UQ>�1Gl����<�z�"k'����i����p%NP���j���dL�RG���[�(�oXֳ�����`�6�>��V�l*m����D��J7��2�ye
X6:L	��J;=-�b��E�'����}�t�/M F����2��z�8'�Y1w5+�\����F�|G�N�"ҩB��f*�o ��P?�/�,;y@����Vڡx�V�.�]�ZY�G���^�#P�F�pL�$oI�;Mq� eɚ>6�s�跞���B?D����@\	����P��V�Bօ;&
��8|�T�?.r��o�j�m���4N�&��R��νHO� �
7��*X�lN=�
<���'�z�
�^��$w��Sˋ��D]ڼ��P��?�,Gm�;�0��-� ;��(<Ѩ�aL�J[���^��᫳*"z'�9am�.<i��l�o&x�;s@��{X-�6G,h�}w���d���Y�O�(D��fd��v-��1����!'}�P�ۂ�2W���s4�C+"PB��Y_�`i_"}Tv5I�@<���=J%��b^F`�R��dQr�Ĭ�U��^�5�r��]IW�S���v�I��{�� &��8����v�*cD��00� T(��X>@a3�v4#���KU�<��/u�����i4��"�3&��Dm���[i�g�ތ��G��3��i0
��7L�)�М���y�!��\��Z]i��b�����v׎��ܶ���C}X�:�^N�&3�@��uawyƅ�M�*��(w�]2��YTP$+��cΖ������\������]���	V@9t���eĿ���I%�RD!���>҃����?���V��>T���vT�R����0t���#��aj��X-b��8C��X�<W�}�n� A>+�Ysj��m�Uz��$ҡa�a����l��vh`з�����X�K���u�W6
&���y���M1x�.
�� (iQh8����D%i�lxi�L�n��6qy�n��^o�<�a�qA%	�
`�e~�����:�BN�K�NP4�����^�>�EӾR�ajL�s�����S4q�Bs�&�~�g��^�<�K�T���s�/�r�����aQ��0��3M�Y�^�e;��F��v[�^���Ox���q�s�l�}�4W�/�>0�p�d����2�@r���vO(4�
�|%�mdm\�;���Ck&�z��K�55�w��]�5�AP��`���7 ަ��E.�)y%Z����Q�Ʉ]oH�h%�D<3ŉU3��<O:��C�h���3�.aJw��z�s�����<٣DpLQ}���B�k٨���+W��������y�.� �q���<)�a+�y�dC�S#V�l8� �i��To9:N	l_���_�����4S� Q������1f��ex��%ۭ	��{�IXN/��1�q�"U�E�e��˚yc"�uZJ9'h��a���x3��۔�aG�L� ��ױբ�1�[Է;D���;*C��2�WUk-fM�#U��'��:H��w:�5��29���z�%�(����dSݦ��%�%z��n��� ���6�n�dufL�	�X�?gl�O��V3E?[������4/3��:<0,�l�ʞ�/�@�NP�I�-ul�L^��=dS�Z1�to"/��)����:G1��	&Yd?��bGA����8!z)
�Ue�8�%�9#��^��Qu���Q)����/~��	A!�DN�W�bk-.�[ΑX���j�&���h�E*Ќ�W��ѦG�ĵd�	���%B�D(�O�����r\�����I��%�K�RF�*�m��b��.,h�i��MJD
4�䎴V'�mp�=<b��wP�Jw����?�l1�ķ����3�?d�9kaT
	յ~P W�ɶ�ȓ d�� It������.I��3y&2"�v2�]g������M9�L��q�!=P��8bK��O.�����d�C^�o�60� ']�P��W�WI3ީҐ�mg ^��J��[�r�3ڽ��kd(��o|�$��}%F[�1��:'��^�$S:���}��@�^Y���������&�x桅��r�T��	mDI�J������nhiw��	���9ίJe�x��ퟺ��p^F6l�b��beS '�щ������?Y,�M�4���j��
00�v5�p1�����R�։�������ҥ���@�s�Tzi6�g��b��+���ήf��;��$-,�c*�޻,�]��v��%����B�h;�c��lp��ݗ t�z�R��k����Ab4Y��I	d_��^ﰱ���F�
�n���	�8������.!��g_I��\�Z���2� ���)Cwō�*\G�.)�ֻ��k���o�GF�D:Y��ը���Ȩ�BNm��Qye���)ۯ��U�P�%қ���u���-a�,�2J.�1�:��p�m�K萲�x��F\?|��L���j"����"��6Ľ7���皎��_��}[��t��M<ν$u�����ZnrHY�/=F�k"b{%QF�&\�y���Ɉt���+�a�^���"�@���כ���vX<�����<�����K;d�@�oY��<i�W((!��$���6��I"l�b�?��g��j1��\F�"��$~�#���O=K�5�ѽ%kV�iޟ��Y����z�ϫBE�jO|��$���X�S\OM6�^�Ĺ���?����r��4��_���RK�� OO3PB�d� �|m��~��#��#(IP���ܯq�FfB��'�l�cAf��)�_�9�2�Пi���6��YZ�@�g�������+�ӕwj�'�h�7\��;�3��Cv�+)f)��TBP	R���$ϭ2�t�MUV`�#�+	��)�T���/�ȹt.?,h�L�p�Z�A�L�'Dǝ�}c���+��j�*�w�DH�Z{R3�_�Tl��o���ʡ]Y_,�5E�~E,3�2���������n7W�Dw�/�0謾��"t,8B�S;��m�z�ys�M^)�5�E��M�4�/S��^<8a���pE�Z�֭.%�ac�;:�U�
���C�ZYH��Q�Rp�i^��H�1Z����֖.u���C�ˮ_Y�ב��f�+m<[���Ԇ��lk��u��K�$(��Ї�M�		�����Z��d�@2��W�TYt�W
FhxΘ�8�Ui��#����؎շZ���i�-�1D����sZ1ąm&46�g(�WkiWU��hA�N�}��x}��@���cD�����j~�].��vzL�5y�礪 ��Ǘ��H[ۀ�o�pFYG˶ėrn:^�lY&���Oj��?��!N�t�[��N����p��w�������K��]��D>�!��#jX�&���V!w�����\$�Tm���B�U�G��D�|q�k�C�j-J�%-m�W�#�k��~���H�_Q19�-�%Z9.0~�G�YQ��*8ME\��"����Q��b�C�I�q���+�Ͷkt:�ǿ���c	S��� �_���#�'�Y�B���Q<_�.IihƼZ:�i4O�E�-�-�okp��[A�/a���)~X���z�7����^�^{?����V`E2-�ۣ	�C�����,���ղв�#���+��� ����Mf�\��a�o�{�F9[Uir�4�Md�����A��*���\ӱ'FB�2�_�S�z��PF�&�O�������g8�L&��"T<���Ys��9�P$D���ANf���bk�Y��6�l�e�;�Qz+�Q;�4���@��0y��G�\V۠�JK����݉ɻ���Բr�&L{/R}K��b����T�ԕ��"�l���?2�N�>�(�������|�汉M0�D�\<���HF����*������C��'�y?�3�ѴQ�ho�㵁�n"J� ���W�����T��=�꙼��a�}�s��ى�e6���ӕ�$l����Nh&وF�fz����L%&k��6?�sgHg�	9˴��WE0�l����t��/=��A��i��n��y�dB��1i�(�9�����Fq�Z����zӾ���!W���w݆D�3nA�,�
�R�n��^��\k��t�1n2(�r-�����Roqy�R�gO�mk�!�N�Qn��n�ٳe�_�<�
5�T�������=P�'^��(k_�m�l�ƐU�� �
S��i\Yt���K�&�L�:v�/�B�4k��}��a������L��B�R׺�q�B���n�J��џrŠj]ؒ�k�g�r����*��ﶡڶ1��+\�@�����*�V��.A��f(E����f�BB�DA�{i	��f(	�zh�A�繾���̟9��^{����O��wt��И*�wT~���?%)ģ�<��m����o�&s�_p�:w��"���)����Uq�|��'�;����Lm;�ģg}��g�t������(��3�+�P̞����9IX�8���t�![��r���/BK���U̥B�0�!�����/�_�k���l�zVZ����=�Ŗ�NV�I퍊\Nò���H�,�;>{�(�������\�����˜S�?|9���ч���lR��lz|��TWd�'���SF��E��$�N�`��w�X�ٲ��h�ڼ������[G�o�U-���	���p����b&��	��������է��X���@YC86��o9�=rټV{�'%�Е���Gw��'V-ƃO%wU�z�c$�~��?Ir�4��>����<��&�:T� n��&�Y��~h�'m�ѡ�_����8n*7����B�ê����2w�E�J�3?���e6m��Ӈ��f�N�X��ֹ��~�a�p�:��%�<�%]�D2��gb�2���I�(�[�O�o-A�m���=������ܻ�2�2���UR��?��{�I�<b]f�43+|��2�@h	�q˽��uV�!k����2���G�+N�{i�I��s�w8	:T�Z�#���r@q4y�u+���Ƅߵ>�SWu��䌜�n����t�I�;�vX�U+�ǂv�q-�agQ�L9|O�c���_ͱ�t��Q��)����F�-1��U�ڴ<�s�$T^SO1�K���&Fu��&��6��|W�}�P2�D9{V��,�f���߇w�2�2�C*�p׳^w%���,���P sUw�.);���)j�4~�t��T@Xk���Fm��0�b�����S��q�3.�ذ�M䧅�%1���"���eݾ
�T�籇���n��_��ȚR!$h��xD�lZX�	t��7L�oӬ�:�>����U��������@�՚�x�=o����ۀA�f�ӌ��C,FZ�Le��?��["\V'��	��uS�3ȔI�RS����I�ՑO	}����ɑ���³�0����C�r�%C�Ig�-[p�˵��O��)�_����U�uݪ%��
��HT�Y96|g���Ǖl�����XR%���QhA�gL�T�$D�@T�MۍȊ���=DM6�~2���/�X�Y`ʊ��	��!w)΢�[1�u��NU��I/6_�қITY׈�8��ÚT��N�ea�u�ę/�����̀��$�sF���5�)���T6���w���#������z�z<R��#�*J��靸�ǜ�����|;�6��L�_Z�YL��@26̔կw��������S{(s�žT]��{���>�j���d��D�������/�u���p{+�)��w��jn���P�^���V�������<�M����
� ���]bskQ�4Ro����u��Y��A�aj���л�5�]∇�{�FB�+1_��pp�c�c'/,�+�o	&u��^���Yʻ@=��F0<Et��J��YYI��|c��S]K3o�:��	|��֎
���ur��X�9�D0�ԃ�K���-�/q���,-�A�z�6HA
�I ����$8K�� n�n�rleI��}��_,k��U��J"�6�х>��S�a��?�)��B=�J�zVNY��cf��5��v��3�b?��Cc#ļ0HqI��L�Y�vE�N����3���ݗR��uɁ�?j&��Q]T��,^�r���v|%�\�>�о�!z���7�*�%n�gn��|�'�J(�ɛ#2���#k�{i��$p�\�ȅ���X�@�T'����l��O霈��YڰJ)��H�bOBU|��^���d�<S�vZ�K �m�q�A��u�`����C{�s^��H���N".o���b�	���+y>2o!�٦��~C���Hl��K��:;�LU�Y�[��yg�귎�;DsPM�n��D���#/��/��ۍ��=.�����?�)3S�7�3I�����k�j�xP��W�}��i�;�#��{�]�D���+�Y$���6�GWa�z���
+�����z�Ё��߹ߊ�X���_�ˌ�����f��UT҉5;T��f?RmJi�kx��/@d�r��Z�"r�z�)�U�Q�o���M_O�޲�Gk��8�^���q�C��.`oeŗ	�R3A�%'̫��d�IU�����[���ɚ���S�A�9l1*÷�Ҋ8ف�{tf���*���n���q~�:k���

H���4�&i�4�׭�~�5��-�z���.���60�'������w�45B�
�n��C{	 ���������So8��n���e9��������O�5և�ǣ3ر��7�����[��	��K���;�*�q5	�\z�j
�3��R�8��Wh]DzM�����"���8Lc�����@U����^,C:,8���$��N��*)G�j�.�4|v� �N-?�r��5r��l���[M@�E�'{[��ɾ�U�@�G��8����E���G��8���G��YQQ�� ܛB
M�/�d��V
���=d�%?
jYw|AQ�->�R��ƏU����^�Y��g|��Σx܌Zޭ�и�؟+�t@�K������m�Z|�]�
��H)����:�\�B��������v�]\k�����iʆ���-�:.kT��YX�m��*��0g���$M����2�T+��S^�&���w@��L���K9��bV��w_�j�AthH��
��uȨ/?S�S�������Ϭo�ǃsk��(�1�-�X�:�p�4/��9�<?�R�j�AD����`yS,˘}���8:����%��>���(�#�fV��).�������nN�8-D�$܏O��H����+���E4��>"�5���0V�|�r����/ٲֹ��+���a�IE98#Ut]�f�2ܣ,�ʻ��ړ)����5����0�����`*2_�`7C�]m<e���F�µ��}�p� T�y�O�1U��:ݑp?�[�_e���{�շ��M�}m<"�NG�>��I��6\�c��� �
�]r� ��e�����iE�Ʀ�gJUiEnj��R��0?��  ��ef������jK���I��#$������p� ;��X~&@8˜�1#J�fMÀȱ�V�t��	��(g�XY#����7�g�E�9ծֲ�Ψ&�����=�u̲��SNK��Y��Eɸ���R���+��M�c�z�,}�zY�W�Cy->�l�Ya��AK��"O�̦8U���X�>�Qm�%�m�<� �x�?H�]f�3O ��d��hr� Ex�]��*��Ƃr�Q�۹+ �K1�'��&=K&6���l�O!����������]��]��s't�<\�5���q�^EXҖ�)���<⧼ �	T���~��.: �q�I����S�C�ڊ�_Ǽ��ʆ�ѓ7�ZsT�'�.�3	��	�&E�rE�o�nfPl��5�c��uVz��(kR�W�t��ɡm�qIx|�q	�������=x����5D�~ sAiU��b����Q��JC��J�[f�ZAx���|�	�+$l�dW�/f�����!.��5��ˎ�~�W�0����6[/>�]�{d�7]Q}l�ܺ�1����{��Զ�Z�ﭻZ9�yAݾ�F-0������!���:����t�oZ8����������Fi4L��~��:a���Jv/�Ip��UEҌ��;�7kگ�B��m�=mV����Z����k36��W�	oXg��i��?��%�b�
�i�bf�t�1h�C����ަ�uܳ�������ț� ?ǲzV�o\eǩ���ٛ䀠��:~~�����k�&=8B���E�ԩ�=K�SwUJ{��7
=:�������5M���I˛ym~�w���f
;̬W�l��}8$-Z����N=����?秘�Y����V���_'j��C��8����ZM5���#}��z��oa�r�W<�r3<<�����eHxp�8�>:�o����z�^F�7��E��}�2bbb[����V�����m��~��G�}�":�^��թ�杪��"HZ�4V�4��'>����n;L����:����!55�]�M����:eK�szr��;��B��a�a�m�O�@HC�]��0��b�����O��4��L�)I�[k�;����qDh��pD�Tk�_�ߴ�J�,ڊ%������rd�{��pf���z�
"��5�&o �AS�/bߘ=㖙b~���bs�`�6w�i;fi����(���߽u0+xC��
}��Q�a�R�J84+��A��.<���z1��c�ώ�>��Q�x�<|�a^#�h��6�w,���y��@#��yF,~�<�QʿL]�?a��c�;и71���"�20Z�K ł/�q��,}�W���Xh�{��?	�*(X�Zp��so��#wN���ޤk�)\�!$inl|ӝ�o�����`�ֳ@/��y�>�q�'�������݈�O|���	�4�<�X�A�u	p�"���O�x���k��1 �)#0�{��a$�z���e�U���D�,)ÿ�2z������)Q���7�"�?����f��\���>�ٞ�^�sQY�>���ӕk�]���R[M�a��WNT1��$0�U/qF��8ٰ�.��b�HA�A��_�jVv���<n,czP/µ�����(K�s�/�����V'�P�nڋ|��}<F֞�ڵ���og�P޶K�g$Yo����6,.U�w����	h�pcf�ψ��,���I�b�_�>m����ʻg�PC3O����7�{,c'c/�MbSa���ċ6��{c���Ɔ�Y+%�"�i}iR�X�z[yŻƟ���a>��)�iD���9�^w�[�8QIg�ŧ'F��Ws��Y��],�bB�cHF��b��/���|M��g�S�Svs��M:n&* �7��t˱��fS|���~LQtho�Y`Q$!����a�2YN��'�(v/"]-��]�0nW���_��b�@ب�����*��"�zNuU�մ�g`��:6�7���'U%����م~�zP�[voG�x�l�_�U��R3=��� '�ki�1%�Y����:rꋾ'��}8�	ˊ;��шE���Pس?���7��3x���I���>���y���tQ��"��K� ~�.1��4���5J���?��³����J�`$lvil���"B�ǳ�Om�-b��ʁ�ZIY���y���Vn�����i��;o;��=�z�t��u�d;6�I�-zj����M�݁�@�7�<A�^����o�E�U��baY���#_Bmj}S�R���u��Z6����7NW���z���b2k��B^M�����_�k�PP�A�Db|�19�A\�E��J�n�Ix�W4�/>C~�-	9�_�Jɔ�X�B�MѸ�=+�����t�u�������z���4�-�{p�ML���G�,'Ye����[��K��|�$�={Z��%�ny��hY����R2?K\r@�7U�����E��ƐE���
�t|q�����p���O�*z���0��z�Tt���@X��%��'rߤ;��[��5�y���^���=������l3�W���5�̓_�8�w6��/C$�yE����;k,BX��e�|��0�X<�T|�>�?�	�x��I�Q%���7j8���|�m��K��5������c��WG;VY�AIͥ��j�Lש�q��,3iM�SA�a^#��R�UJ_�4Q���7��K�b\�Oc���>L�����g���'(�H5f���W�)d�߄�w�ȵ��7�Z��B������f��0��`4�ܕ������;�([U�=��<�1����l���3]���g{�5�F�i���oթ���g<N��X��P�%���.���A��b��hвq�,���?��Ԭw�j���n5�ԑ�+�\�>?����|�u�t�J����U��G}.�N� `yZ��O�Q��~S�}�g��dF��`�4�Eg��Z��Iډ,�,�U*� ͫ<5X�A4P��>|) �|���>/����R~d�eDC��@ͬ{(�
�>�ZT�.º֞��-.��ao�m@3�����0��X�@w�7Ҭ���`���5:�y�N^"f̼�V���Xȹ���p�[���x������΋-!#wa�e}���]�>�z�iÐ�N�n��1�t��"%��~��u�wb�̫���r��5�7�Z���Q(����%CCjum�����Z�h9	��AGR�Whp��u�2�8B|γb�o<���,��7y�0�� �a 4�d')�;�u�J�����r�[���8�v�Ƙ�l&���=L�R��!#Ѡ��O���Gm�ҺN�����%L��Z�RoYo��r�\����(U��kk���Q0��=4Vv��D�U��0/�!RN>3NJY�h�2-]���i�����W��0V�<�a����7j5��&"��R��j�)��s6��=��~{9����8R�A���e�ݘ��Le�N���0�C��&D4۟:���e�D�ay��Dk)(�X�gj*�Vz�ů�f�t(/~#8j��C�'�E	)��2�M+�ҭ��x��z������֣;�����*�H�V�J���4�~ 渘����w��9����R��h���Z�F��&,cdc;
��Pl��2��\H=�#��i�A�`~/ ��s�|����Se=w������v����[�J�.�č�}HI�tKj��Z����2I�p��ZvW�TN]�n�Ā����/�̛9m�؉D�XՔL9�<�o�0���:uN�}�U7�i���',Pl�_MM,SU��)Z����y@��\��/����"y�-���(���y�P�~́yu� �R<�ԀO@�u�a9沦#��Td>��{ݳST�8����>/�S/,�>ƫ�"���٘!�4��
��4���p��>En�bP�B,�у=��g|�*�9ۋ��&��/�B:����:m|�C2d���l��i9؍��	G���_�<���b��փ����1���i�P��%�ǥs��;�q�M��*�K�4�5�֒ͺZ�Cɻ�}�����Y=u��8{g4�)��~�e�mVf�g��Ҙ�Uf�(��}h�^R)�����M&G�$��m����=�ܨ�{��bT�O&�w���t�ޫ���!��÷3[�X9����E� 2��z4�s���.7��4?o��+o&�7*�8dF��+c?��I�}���A.u��p���������{�?8�È���疠?�7��f{<W���9�5��*b�i�WQ�������o�!K�V����`��
x����G0������vd���楶b"J��]���J26�A92½���C7����n6�d6Ms��)@ZK$C�ᕈ^��5�w"γi��ח�1x7_ '�ZOa�y�}+3�!���7v��r�	���=�$e���e}l=$�?�Y�����\�=��l���zf_��*b-�6�Q��q�Ѻ�n�9�2b���Lc����礓
W�F�c�$�9l�
u|�.��]R{��q|W"/)���}���.T	ٳ��#�T\��1x�4='��w�AG:{'RW-Z@�v +�j5����x���2��l��e��Y�; �bnrHu�Uv���i�
��<v;;;s���18�M2;�[�{|��2%/�U�C���-�
H��f�.�M�'.8WE�uQ7��o��2C9��gIm�~|kj�԰I�hg�75�Yyxŗ�c�*g�nw��}�9m���Y����83OXG��008� �푴A���~PY�C=�u�����_�#5�yp�}�I�� ��w ��O{�����r�_��!�hʯ�l�-����qoڪHp�"zt�̴�6Mr�e�D���2J�I�	�N����j?*���� (����a��?/�d�$�3g�02�Z��b��?��mJq�}����^����#��c2��P�h�u�qq����oE��a���W"j���ǑI��-U��K�[��O��	�ond�O�&29F	�w'ܴ
�%#�+�^���ӜIi��Ȟg�~�f	��M�T�~뗩��{ g�I>�@-�B�X�߀���o�ا�븿�n?�0L`����yϠ!���q�,P될q���3Q �����F�p߈қdK��.xNA���U�aY�Ӊ�7��w�䯫C�����i
��� u&!+�1�i�F��k�Mv �[�:�IbTT������$���ƧjV%����s��aJ��0ޢ��T��"�X�J����]�k���ˑ��b��+��=j-�,;m3���-#��[�*BS�4E�L��J�n=?��p�l�����o�����p�^d�j��
ӏ�b+kk>��'9�;�
8T	��~���2�-wT���46�p�y��4�ֆa�U�6>Rs� ��y�L���F�K��}TF�c��*��$4�_���s5m]���R��c
�>�E��: �J!�:���t�2���4�.�[��mlX�.�giߞ=-G1���6�-�U�Zco/K�+�o2H%2d���u���}����eӥ�i�%���e�H�U�<m�Ư��S��ъJ�f�ce^�?��8��t^��p��0���n$�}`ո�ʣ�T�5 Bd��:�ף���
�{7y�i'��@u��)��X�	�Z�u{�й���F�ۆ����ޡ�̿6�1X�k�KH�JH�N]�<VId~�
�
�2VϾ[�h�?��g򑼅�{yF�L��D�'d`iŀ[M�n&G�#k)�e�K������f�/��=�=�d���3��>�%X����
~f晋]�ӊҲGS����~A�H���<1�I� A����������BDB��k��%*���]Լ�[7�Q��X�i ��whi�g������g�0�C���"��]�f���2���*>ˇߌ�y��.I�T��f,�U����Oߎ�Z�W1�06�\n(e��셔R��du��1N�嶫���h���G}��X��w��q�����~�l��� {���l�5[��ہDv�Az�OnZ�f���;��W�
D���ׯ�"�2O��)~*��3�U@���|����KK��I��È��
lʫ� ��	�S��h�+�Q�X�h���$!A��&� 0��3��vY���=rN:����u+:*wY�����Q�~�I�KxE�EdݑN�ܯ���>!������#�+�q����&��oԹ�T/��1�w�����_�Ft�D^����2Y�����6�9j����%hRH	Rތh��A�/�`ۛ�ra��ZG�����=г��ExM<�y��=\����؇��%�$��w�N��d�u���ۄ{PN��b���+����Ne���
�x�{��r����}]���Ayd��?�sh�������L�\1�yL��[Sz�G��&=`���׸t,;��fɄ-�M���۩<�K�^�#Veggۉ����o��#��u��S�S�B���� 0|�W�#�ۗ���~�&�+*$��ZLj9�:4�8�!G�T�S��7ٟmB&�L
�Ǆ��8���M���RE����}]�R�lW�߮<+>"�>�yX�yd!��X���
?�c�������s�e�R��rX��Q�s��9��3w��)�E&�aQqp?���� �5#omMG4���E+���%�?D��x&0}M�d?�h6G9��
�I��%'2�j$0aHj����W�t�ϓ��0���:!|���Ԕ*Y��g>h5?�̦���Ŧ'
�:Q�εg'�"�_�,0�[�@��\>\v=�,ϑcǅ@�chB��a&X	���O�]>Թ�QK˸*V�c)Z{4�-ځ�?b�m����6���tE�BD$)�_
�hmOMi�H�1���7^�+@��Ƣ���'+yv[���$�_^�&Z���n�ݑ;/B%`�%��}��UZ��ZN��k��k�Є!k�u������Ac�9�z;EÚXD]� �}�͢����Ï����GD>��]<���-f���m(�-�)o��?��t�����C���|�34O}K23^��D�;&b�v���T��E�M�����Nf��D"�K�o�-�;k���F5C^��蠲N�2�^�8�U�H6�f�����y0K���ڰ
/թMG܁�z��&����[���d[����)����.�6Vb���AxG��YKl�W~��wH5 6��h�D�L��jV>=��( ,�z��o�MR�`i�Y�[����ad��j�HS���M2b��[�xg����Y����3)F�t����eN�ZK�%�~ �w3v�eC��?�ʞ��&�\^O؇�x�r�:X��XK��u��a���3������[ʀ �jM��K�q��F+D����|iAQn㡲�ڽw�����ɓ#�1�/Mg�O<�;Ӟ��36�c���#�߻~��_��k�s�y�ʶ7~��L��u�w�T���Tt���s��%:�Q�M=��=���Ԏ�Q�H�9��� �'�\Ȣ���Q�p@���� �_o�H�n�/"b����v��*�5��>�f��S�k�V��y�:�W-�R��_�AY��qxxxZ�(�Q�Ry�������A^�����
G�[����73�3�#���7���N�5!j�z�r�󧟣�\ K�^�eo,ӼsЙ����3R�|j��j> �uW����N�`r�+s�*�Pur���#��*1�h�]��+ a;@ݝ����7�8��h�!d'�E�@\���l���On`��^>��K�42D�z��=T 3���l·">,&�Z����&b����a�#���o��J�ť�d�\J2Uq�f��jL��3-���Xz�Q��2�[��<�C�Y����Σ�*z����ۓJ11~/1�ꌛ�r�Z� Ֆhf��*4e�h�P��Ɓu�/��C�f�B�?��o���Z|� �m��M�^��)�7ɗWuum��~9���˻��֡��vl�<l[��$�S�e�+ü4�z�ś2颕�^l�.� �U�
*C��g�9:��jh��yB_��;(����7�CP��M(s*��;� �5���L`}ZќM��|��[��4�
�����* ����_�i���/�ͯ�ٺ�a��o�~[g�(�dP��Ö��m���6�0���xc��_e�Z���|��ј��C��X�4�FJƄ�:I���S[�\�z�˝�_�����}UqAՇTtF�V�l�AF�;(V���4�uǒWP�b&�&ɡ��c�V�4����{�� m3H�VW��*�ÂR�z���VX��� ��k��׊&=�"�|4r��ׇӏ:���3�$,�N�@���#e�����W��y�s������Ҝ���q�0��<%epz���+�߈]D�\�OqU�X��3��a�QE>�+���ER}�J��9���R��B��G����c0���b|�GqV�z��]�X.�0��8��Z���U�1�o��+�˃�i��ʷ��@�����Y�㖐�o,ٰ�_"����<ǣ���*�M���,��i��	EqQ�H@WH����{X��ƓO����P�U�uum֡�ݝw� *+I��9Ľ/��A���I���i��s�v�G����Ɇ���_y���.�x�9t��\�#BV�|I��R2�������!/�7�j��G����ΠoL���������8�:�%�4 ���LH�۴��SDM,���+5ni�-��8����/(A��5����,f�3ʤ�ʪ�v�����p-��喱Yl�?��X�C�;sV���N������l�] \���&أ {(��s��j�Z�ϴYzݠ���CV�D`.�Ğ��'��8��}������$�c+�F���~�����~סwU�F�w�iC��\>Eq Qד�9+��}Yh%3�/�U��^Y�Pr'�������c��:�;*�\�0n��@�d�'�t���++b}]�?J���[���j��(YԄ���k[�w���E���%H����I~��/�������ͺ숙~�d�﨏��L�d�%6%��/�*d1'u.9�|�aFS�����)��YA����d�? ���>W�)E����t��x�~?ow���#ɳ�VÊa�`��B�������>��6�9$I;������?�뮭�����Le%wq`J�~�d�E�v�-��JN>0>�Y�W�r�[��X�~O����"����l�5#G�83k�{
�Ӣܛf�%L�?q�|����~���)<T�N�J��PG��Ki3�����!�/� �[���D3ؖ#�}HL�3�᛽X�����Q[�n_|��O��!�>�v�9�ilSb�����@��y�-fI�33l�wG�;�j�����s�?6��;�bV1��#���y(ՇRfU+LJ'^"�B��vk������B�	�$x1�uy(j�`����nce�m���a�Cf��l�ڿ���2vӠ��Zm7Z��H_qZ�P���د���3$�v.���.�SU����;�ĐrD$}cٷ&P���y*x�Lw!��rlHL��a�8��>�tM;V��͍��D��W�c'ݙ�<)�>N�jk*���%G�8�4��wR��w	l!���`dR�AW��$ʿ-&��f����2B�������o��.�����_uG���o`YC�M5=��$�z�H�.bS�sC��e��/�Ї�Q��+��+�wD����l�k����'0��C���\!��P�)v�{Һ��u�S���,�>F���}�B�� 륧k�$B +�-E������>�j�A����>Þ��a[~�����ǅ�����]s��~�5�3�UpY�xw�6�	M]o>rh�kV���:w����pu�l���Hxe"oؗe1%��P'U~��4� �
��g*�&���c��3�b%`O3��'��y~��TOl5{3���wm�s񀟯$d��*���6��*��Dx@UW�*�P}�5<�)[��1����Ow��u�]�LH8ӝ��!j�%�_��ܗ�2�`՝���tԀiv]�C6%d�K�Շ�H��zt�w���Q����7�e^�.^[\d�пEZ5�<j�����IV)�ʊ�����$�<D�-��_lB��/3{��"�0��bp"ry2+��A'���K\� �jNy��:�H+:��蔳EQ�[���T��q�n1s��rx3�\��W���o���R3`��^�~r�O��5�j�H���Wj��w_����?t{0Jh�A��+Xh��L��`1}j	��5z���'�A���#�c�d*� 'A�\�f���#b���JKP���Z��9�վ���'Z�^�/.�98�r^md������2�x�.�n�φ�������YG�G�������'�)@9�����/�@)洆�D�)*�CB<��O�d��H���	�5��ʀR'|��uZ�%^q�W��N�X��n�ⅨXt/Cg�bݢVp�[Y^t�+m�A U����1MF��&O�3��-R��Ӽt7����d�4��aZ]���U�Ȧ�B�c���{�Veo�a�H��J\ȣ����oRk��s%e�[qi�%|'�;+�3_rX�
"vGNW���|��7&%���ߤ��k=11����m��:#�������?ox�+8�/}�c�}ߒ�튉����\�*��A힇چ�s�033HW�?�%F�UZ�k��R2�t����CC�({e������e	 �}�s�Gwj�S�f<�ƭ�$~��O��]��J���B�"�ɷW�O�ϮAM��i"�sv���"�yS,��=r��s,�L{�5,*� �p�  �L^8�ԓ���,B����*_�7�4��/�3����42M|���8�8'�+9�6�%�λ�/�z�k`�7���]��J;|�S�5���A�m���������u��iR��,P�&��zR*�%"���B�kfjI[����c�'����B���<A�T�°��${ǩ#s��ܞG���3�U����1w�L�x�\��B5"�mV/G�]^�z�2����o��|�g�����si����?��z^{�B�%z��]5�+��/�iXZ�T4H&�ht���ڣ |�Y��x���,���0PG;���0r��i��2�^��l��x�Jv+�O��N)����T���<��FP`��%�o�!��&���Am��ky�%�߻l+�8H�l�
�/��Uz@c,�ư5!�8���52ɣ�����UEX��ӷ9�˭�,��M p~�4i+tకU�-]#�l)�GYQG7���Uo�>}Q 5��M9�B<�J�0�d�w�8��Ȩp4�:`x�:��j#���^�A�5��Zxe�IďjM��s�ƹ�=����x�1C���"j��dk�oӆ�j��S�������^����l?��-5B�yW����KG�5)R��r�`��XxAԜ���	�����wrN? ��YI2�����L3[�r6��V�u�?^��A�a-���R)i{2pS���f���~D�~%���
��(?V�s���wS+�����_vU���c���T.)W�q��`
)��oը���ϯA��s|�Dt
AU����%@E�J�,���U�^��39�t�HT����v��<��<؝>TD��-輄�m}��Lu=+�]�l��T�
�ɡL$�u)#EZ֎*&a ��� ���?��&�'��X���D���g�j�%��o��	_%J����D667� �� �];�=��ڜ
����/���E��VÞ�y��i���~��	�u��MлFz����W�4O�.O���eӬJ���9��b{�/hxfh��)����wp =s��c��Q���n�v�a'��)!L!����ϗ�,���Pwi��6_�dD�)�5 ?����p�X��b�R��|���!q3`o�ޅ����� ��]P������ya�X�p ������SI����u)|�c_�(�7�#������O���
��zz��(���P5(�X1�.�bU$¡'T�-�;�FE2ь�NM�$���>�UV�w"��[<s}���d�=��rW����޽�Ks��V��D��{ܕ{7�h" �ń���{%���^�r�i��>���0�Hr�JM�(�[4�\<��'�-=���=�&��h��l��aLs"���?�k��~1 z����m�*l�a1���?�醙=���n�N[�k�Y�e�"�x�U2~���O������A,��G���x;��nU�����Z��˝�峒��)�e%�l1Zܛ�Ȁ���i~7I�T�2�z7"�-� ���C�
��_蕼_�����0hU��jv�� �������g�t�Ǥ#P��󿷋(dǌ�\��rU_�P�J:�qD����'�<��H�U���%�]�TUN�`='�T� �=��0�
�K���c��6e��Q��'�N�+�J�!�c~����/�1�rd،p^���"��&�i��pcƐ�ꧡ���K􈾟=��{�@�`�Z���N��,x��������p��%������̻wr��ܹZQ����� �f��aU�K��jcL3@�̟, �U0��L�k���>�YĆgTH�w����*K�p�n�=�4$E��P�㷺l[UxFtlp 8WA���Y��-��g<e��yNd����$k��Y�ӈ𻆉�(��͡|�����v���"��ѽf������
���'ݖ[�'�I/�oз��wV�s�0��u�k�ul=Z�r�u̒���	�K�O������{�z������m޻�,���j^/���3�<�}�Y�OC�ugm�A*D3�8����q�c*kz�Я��V��r���lR�{�k���/�sa�+6�t��8ӎ���ƔR=o���o�)�0W'��q�!��<�ז�-�8�,�����;�|��P�l�g��K�❱�1]h�4ԻP�yK����>�[��/3�������Mw��I�l�D�>s������mp�޳�59������r]5uuKGG�TU���|>T�U2��ꢟ>�Ud�2Φ�����Z��l�
=�K��T�4�Э�p���x8T�w�b�&���D�\��4#B]8�Ӧ%��y�A�s5.i�n&�>mU'���5��j���'ٓ>[���j��C�{\�d���a�����#��N^AW�nvv�:��Ƥ�ώp�Ʉ�s�V\�櫛�\ѹ�w�[���_s;���Ͷ�����!��N��W�P��eb H��R�K�dd�.�T�ȕ6�Ȗjk���ՙr]z���;u��r�	�&`6��s���ɔ+Gz9?�oc���L�h6��5�W�iu���1�t�Q�:2��'��:s��>��a���r+��9�OBU�n�t��m�,����9[^.�5X��e"I���)5�;��[s=b�g�\�M��L`'��ʚ�bᜂ�~�c'-��Q#M���Cb��el���?G-y�a�E��������'^����QQv�ޤtJ���t# ) � !�"%� Ҩt
HH#��J#��H3C����u�\�,������>g����~�����w��qț����Q;����kO����[�$oo�������K���"�|K�= �$}�52%�nw���;����eec���UϜ�0�;���0�7۵�����A�����,��MT��~��"MJ�Ŵ�ʮ���S7Ѯ��9�˲)Ͽ�l"���#�:����aò�sM��fb�����ô����Pl>~��S8���63H���	������6/�:��S{v�EJZ�.o,Yf��i�#`'��|�QG$J�J�'Xc��\��d5��#���) ��K����Ff>��}� �Jz�7�X3�Gk9[�"_س�E>f��Ń����]f��𴴴\dZ�Vs܏���n>~l��,��a� ���ii���%��@��̖Z���xD�R����*"f�r�b}�-R�8��}��Q�(s�!9�)�۽��ז�8
�Ƣ��.�E��A�������>�2-H`-G�tF��($���w�|Q�tGw��+a�S޳�P˭NP������hL���Ԣ�� ��Ym�Qm4�	&))��������e�qV������#���^���с�Ч �gnVu7��ƫv�O:T)c�Q�n@,��\�fJ�H=<<$A�ÙOC�i���J���g�F���fJ�ah����u&~��x%&_���}d������s�ǣ��e���n�<Z�C�]�<��c�rE��褁��V̧�Q���pU�i��3ㅯ�$��4t�G��� /��uyN��eL�f���6"�OMuup�f�c�K��(d��<OcZ�Dٿt�44;�ҠW�/)�̄3o��T����T�^W��2q���Z�tKv��6�՗s��f}b�@i~pr�����rfaNk�]�f ��2j7ˢ�C|n�+�J%�/�4�e"�+4��-�%Pn�ʆ��7���^;T�jO�trf!_7��q��I�s`�m���ULrQ���|j�Z?F�+�0�-����+��u���[�'�9���?g�m`X�O~���z�9�w����܁9]�����s�*Sh��U���|�s�D6�)1��b�[+��>Z��b7��k5����X�9��o��k�eh���0��Pk�?��D&ઑ�$��ۡ�!�S�mmquuO<�lV��D"�ūm��UU�Oͧ� |Y�#��o�t]�F�ܛ����L���_ m����o��j1F<���+yLo��Jj�'h�_��ԧ����3z��7H�$�F?�]����^<�D=+s��'l��w��(¶S ��"��5��ȡOG$���x�@ȯ`�����>�%_��)O��c��4k�D���I�(U>�
잕�;���X��,�N˿�Z�)&��cҍY?�.P�g+���Cͻ���d����_SO/|��n�c?�tuu��^����>h6���Ԅ��ޡ��u>�WCS3��sn�=�A�Y�Q�^�-^�3vK�����@�Ufʂil�3;�����9�^V�:�N��B�}8��YT>i'��怲��A�!E�x�-&F2�f02�e�/x�
<�7��c�#���u�1�����;���>�Pbt=� �� zSXD�
�1�/��X����67�.\������nF��(��<��HWF��]��ߠ{�3a��@� 􀞞��x�bjj���9�/�y��@�nY�g�St�C�`�@jNN_��4:gL��莎�]W�*L�ြħ_>�)��`~�jÇx�9�����_S��wV�J��d�AZ7��ٞ�*���~���9��b��Kk<���q��M;��(�b��%4Z+�mt��ay�ƶ�gE�������5�N<#r*@�T��.�\1*hZ�L��UiZ>�DYZ.E�l� nĽ��M[�oib�e�ep�,�%�7��[�����M���d|q��_  <<L�-�Z��@7&��� +,Je��g367ﻸ��%�>n����Y�' iMZ|(6GrPp��GF�M"����t��]��h�g����HI���h���:Z#hF����A�G,hAY��/ "�(����f���lŵ�g����׋1�x�,��p^�%�E" ޘ{h_V�;П~k��SnI�F�O��A桄 q�v�n�+8�nL���|�飈�>��w�]u虁�3������66��L�y˞݀&605���q�����z=�1l�A>B��T��1]a�Un��z��O��F�-���#�S6Dx�����W*OВ�2YŃuٖ!b3V5*;�H�}��X?��4�����~�F�ֺ�8d�����}�S��c�ZksZ���<'ǳ.j�l'��˝�J�S���������>�r{��c������^*��r�g��ֺO�6���}"]A���3O���D�f�̓�`�吻^+}�;Nd#:Q!~�h^mF�o{J�k`h�17��I�#]c�/}�X�G)����)��?��]Ox*���x�+�C)��{{{��2�T�"�U�b�S��`�Xꅗ��\̧�;MJ�j�=�o�}>��J�1�_��{�>��*�<pd�,�e���a叝��|��$~U˿���� 	~�����b������`��қpo��^�B��%T��`�=�!"��Oaܟ%��9���Qr�|ի���ᡈ��>�7��m %hii���-'-����X��ֲ$i��o�f�rC�u�K���Zo,}�����|c��t���� ��F��CEQ�FɽI���ū����l��?�y�Z;-CstAA��ј��7Y�Zw�Ozo@��ˣ��C�J�ls~N�ƚ55�2��~��C�rys����;z���@�O�(�ڐ�� r���đ�;�E�9��Z��&i�o��Cȿ������#\gD��a���������r���wAe�k?sO�M���F���1A�t����,�JMH���Nhe���/%��Á�����ttt��<�4n'V�����Gypx8o�é�M��+�N\�z�<6C�J{,����N�A�rV�
�ɓ7y7�Ƙ8	>��*��x/SD����Ҩ�9����$Zܺ���AOi�$����=`�Vf̀Q&E��:7%H^#s���� (X���M�8Qա�;�ڢ����v;��/N����^�&f  �tG����4r�t�����f`b�`j��'���P<����s��t��7s�Е��K�r�I��vO��oZF�LUܲ�c����l$^��_nk�9l�nT,py�:�ȥ{ѝ0����\+ڨ�
p�n�~|i ��hG�e��Q��y�=��WeQ�L���g���۳?~J��}�nnL)��w]�����%�������K��P�w~/�Q�E�cZ�R5��+����^6�{�ō���~h�������$Wpct����Oԛ�����f �	O�1ȀO���� ����INIA� �D7����(n�ۘ�r`�%������H�p��Wfw����i3�+i[�7V8K���F��_�џr����h=�v���	t�l	8�ep�K��COXxE�O�G��m�;a=�@2��F���uV% �~�[��%ߗ>���c=�`VL�2���)���:��R@�A���%�γI��P�/�^>MA�#����m�*����p�V/�}ח(�?�9ܢ�����H��@�q�L)/B��cJ��0t至�}��S���w�s��v�PN��p�q�*X���=t�2�8K��l�Y��H��|���^�^D=�gߓ�����[w�ۥ:��";e���Z�k��j���K��5�z�T�f���N2~gBcsJj]�Oh� T)M�����_pnb\���-ݭ��L��y9�_̅DD��RgȖ��(U�I��9��?�)#7�aNh�$���Q'j)p����Kv{7���R4�E0�[h��<?����:�Y	�u=���voڃ�`�E��������^��MlΣ�~�]��}BV����"��~#�I��%�U��6E�#�s;�q52ɳ���yG��`E�N�����I3.��Rh��8����ӿ��j�u�B���G�<[˷,�z�<���b�;ńz�6����ɴ��2f�徴�ѐ����L�&	���M�s�g(�����bk4��ň�����m����h9aǉ`T��bum^�*���XX�2jE��C�,j�S}8x�z��NAꣃ��W+�?:ۦCͱcIb[M[D[�����&5��j^����|�Y����7���	����򙥚�������b����b+���?���i�d�>��������>\����*��4����1��/ƃ��]s����\�1�����O� 	neoO@DDtv
sAF�_a���S���ښ߲�����Kk ���םD���_O�]��kQcHB�������o��\�>�]�uchb�6v9�r�=���`gh;lv!�Ȟ�i���������.�M�,!M��j$�"��;��l��j��^m�r�v��W�/뙮�����S<i�@���O:9�ϾȪ���Y��6?�9Io��u<ʬ4;���<��I����� �c'��ߗ%���o�<�n�71�ۥ53%���A��pX���ry��xԫ�]���4	{,]W���'�ª6�L��ʼ�
�^�����5���0�@]�87���Ah�ǁHP��5���M:���y�(�v�m(_�.��I-���gE��6�2���w����MЋ��vpg�>4)}����i�MK�S��fg�ox�+��kvN���>�D�ܙ���E��:�����3�U����w|p�S�l�8�7,��\��)�uF�?)DHOQ��N��((���oֱ !��	� ��l�To*���$�ഽ��v��7��-���=Q��Z1�����P��}ޞ���$�Dm�ry���8n�\�Ϣ?��%���{�������Sy��"��*��Ȍ9l�%>=�t�<c ���\ox��:�������S�r+ƪ�>,�zB���g�.G�ss}yvs��4����O�a�ێ6l������4�z�T��>48��oӢ/�옂�`�~��<yA���`�mgC5�;! %!	h����X�G���}�� &G������������e.6lm(-��dI�������^�0��c����uO����tbYe%��.�ٿY�u�N JK���f{d&��!ٹ?A�Tvd{X�_f�M�������/��6��cjhW�||#�)#���`o��-����V3"�55��)���hU�Ԩ�fF�cnݐ�MG�Ю����V�ǩ���?>�=�yJ���5Ɔ.dd@P'Mz�#/3�s�;�������W���=��3��%	b3QOڭOV|��4�^dț�i�"�q�,�������Ht�1Q�y^�M@]ԏ�����M�IK�E���=�M'<�<�	�~Zi����1�gs�L*��� B~ڍ�d���#QMMM��.����=neee��b�;�+�-��5���OK��Ùە
��W����hB�>CJ�wW��
���-�t3]�	������Q�zf���{LWm���ee��}t��}p��'9^�����@�W���N~��g(Dk�j�]�����]��W-7�,��⻊=Z<�����떖������E~�������#������c�LXO���� 0us����=�~KUU���5`7�I�T�rc����;��y��&���m��w������R ���Xy�G#�(��ió4�A���c���x�f1��Q�tKU�^䞴IVM�7� әL���1�K��ǺW�Y=����wa��G�e�I�ʪ�Q�sjm�vn��:uD����I�O1qh�p30�Y\��)C�! LЮ����x����g����	�o1���n9���Y��� ZP���g����Scs(x����"��-&��-�7�u6�����k�h���G�1�ЈH�,��!����s$_}q�}w�Ҕ*?�����^�zD��+J�������@���O���ݲ;�+}(��\�����!~��!���zB�k�Jp�S�o�L���Qd�U���Z�*���=�S��f����L@�W��4�w�_��-�`�����j��Òq�h-�Ǉ�u3,�{Ⱦ�w��r��q����޾I�AO!�M�Jr�%C�D�?���_�-��� ;<�7��%���NH��=]N�����8x���c���ؤ?fXnoq������Qߚ��gU���L5N��7��\����6A'�Qu��x���9�w��F0]��oZ���:Z�̇�U�D
�T�o�(��w[�gp�@��ΰ��9҇
���#���.�'4w�s2e����=2b�-�^S:Y'��/�Jg��7l.�cuɞ�kP
U���s��N[~�:֏�}������1�T�y$�o���_�l[��f�KZ��ze�6�[	~�Sc;R�4h���@�����L�o�R�p��/�`����eHN��;�ݐ�C<w/eCC�ik��Y.�M�6��,�!�Ŋu�J��ٶ؟���G������~H\t*�_Q���ґ��n�R>��!�h�Od�W����^�\��| 9y'N�����F�Zb��U`�i�(�b�Φ�T�������_��my���&|P`�M�P�K�*v善�yź�er��&��9���}`��z�?�!�XhqĶQ�fc ��Лr=<+��U��
����Ϲ��N-�M�+��-�y��/��}�����ѫi���5It7�(' 
г́W�uF��U�q����#�,��L[����e�%���NP�'֖�.���FKԷ�͋2E��O^���z���XI���T���GL΍�&^���yէ/,A�z����ux�eAv�$����{Ƨ���"�~=)ƱE$�/�� ��|�(2&oo�������y~o$[V�%��2�%��A����[DOI�@��8����j�H� !��C�a$Kn-r��-�t`�.Y+�_��� ��������ȘC�;Nv%@!�o(ۯ�11DEE}.��ai���R7oeV���њ��Y�ou���ߵ�v�����Ԇ����o��-����k�5�Z�F��#�����g�[P��{ň5�u��� �v#Ka��L%������њ������r�痊v�	B�.6h
�WK�Q�`�9�-����8�D	6�|���@���_mH�w��Q��2����ƈ����ux��e�E1���K6 A7+7�skq�f�����)o�._^�1ږb�l�4����AK�z�`���0�rn1Q���r��)J=Օ��l=KM��&m��!��b������	$�.I���QXT�1���w�i���V�j��x��B��rR*�'z.��H�9��U@�`lQՐ!8wKWՔ�$cN�+��'�uƨa��ɝ����m�ݚگ�.H@Į}Ք똚�Cgv��C�㱗g[����f���^�1_S�^{]���dw��5W��_��)���#������[��xv��T�-&7VT�Qlz4�]f�vA�J��{Ԯ�G݀];��<q�u3@����!���U����:Me}����C�B�l�����J�!ᛂl����G!*�(�fe#*��{~��U�(�����Ct����� �HH�k��"a�B33�������0��m���ɼ��Cd�gJ:<�kP[n�����.�!e�y���3�!� �}tg�8F����%*��b�����7�zfO�]�cM�>�-���ϩ:-8a���~���CԦn�1�f�*��z������p'?�ۀ�Ҡ���oNѷ2 >�)�zoQ�;�ēT2"J����|���\^b`��Yf��J����7�5:r������*+��+�F�R�t�_a߬0�`��&��|�!1�3���!�,��n����G�o���V���\�{\`hi�k�q�K�!Ѫ����j��:"j3�BT����cv^�.8�H�ǌ������,���$j���[[���������|<r����Cd��ZE�u뽚�`��/���}'�)�a>��s��v�����O���ؖ���U��ꎠ��z����N����b��_���J��"�J�W����m�)�X~��z��a1,��[|Z��-Z~�P�̿9Y��ߪ�Ř���P]�R��������X�3iV���{3���āWk������o�))uW�X��ࠗDd$:꼠��O̬�u=<U׉u�d��Meϛ�&�H��T�2Ƞ� _�ۉ8�MU��*���#�����M�E>��Zܶ����I�5���G����E"�3��c�]��iJ2�o���2?ӟ�\E��ߦ�q1O�x?Auv=�q�U�dUעd�G��\�r��/����M���5i^9^�ݟ��Q�̖ `mq{s��E�o<d��3ݑ����f~H�� �I�����*�sw���9��$�O�x?Ӛ�;�S���pU0�J�q��j����O@rm�$�J�8/m8�����Q�i�|G;#�L���r�� F&����Tw�Ӝ[|����}��lH��
6'k�\�p9ܷ��U� ��O'��c$N��'��Qc=5�(txS%�A�X�E-��`.}Ukn��-���ڪ�)r�~u��C����ׁ�����ؿ�b��x���>-�����KA�����q��.�+�����)��U1��Sm�q)��;�����4;�\��d�a%�Z�O�hꊒ�֗�Lx8(*�qkQ�R�2aΙ�>n��I��ק���*�r��S�����+Vt�b��� ,0�R�s��b��ѱ;3i���+�'�]B���� �F����?�M�W�E!�~������֜�8���,8+=X�P���L����&=M�j�^�
c��I��d�t�[C<w�H��g�僕��[�z�����x����ߋ�����HI���^�v�7To��#\%������SD>�1�5�hee���*w�Cs������?����d:�ު�W%6M��g~��ڢ޹��9�<�8������W�j^\��)8���G+X�����H"��ܶy��B-��rEz�WL�	�,/6��9�R�rM�_��� X�/�^�:n�j����	��7.j:W��w��`~��f��'��[-��������?���������(+4e�8mgV�~GCm~O+�.T�w���a~�%O���G���ˬ�Rߪ�N����3��̇��z����dy��&�k����I��FF��IŜ�)S����)����.ϵQ0����`��f�ă�����?m�}�S�uj"i݋�����؟`"�'D�5�1�$��<:�^�( E����t�d�����b��b�5f��Mt�������t(�P�=X��)���	6�����T�=S�����إ&�
),|lx}�xs�[m�C8����3���C
�Vf��jU�M��[���`�sm��r��b7�*�>�_�EY^���w�7�nj|�Nl{X���N��i!�ǟ�����s��@Q��F�[�f�`�e��b'��L�P',�LS�R#��)�"�����]{V!d� !���_-��+:cF���u���e:��Ԝ�ِB��s��@���'�f�^��J��ճ8?\G��/�/ ޛ���I)�OX������N�����^x�-��G��(��O��@�X�����ß���f-r�o�`�'��<�+����8���W��Y0���u0WT��%��ή8�f�4>WR�������ä,Kه3�ey��F?&��(�JwB�I<g�Ti#_=��Rt�Tx��v$�'�Q��	&��������P]h�����P=��~���?N��I}�X��5̻���J�f�V,r�l�1B��yx,	-$ ��'d��N�$�y�/n���3l�	�M_�M���,�ݼ�B1�W��'����D�.���p���T�C���>���J!�C�v���S��(�Ɍ��7��w�2��u�5&��Z�!?T	���;Bg� A ����[�(?i��Ӣ)����Z����s�:�	h��0�c��~��&���zc�<ztn�C<zi�����c��h*��3�'���/:x���T؅D'�F��Oʹ���E��^E�,N��*=�F��p��k���^�.2�݁�V³(��oS�ܶ���A1!wi����1�=c��x�j�:�C�Z��x�^��������9a=x����A���X��^7���#g
����0=�	�H^Ϲ���ִ�SN�M"�����G3*�Ot�L���E���!�x��������S�z*�A�bl@��a�-gb(Ѭ8�Lp��ޠi#=��B����_Qe�3���#��,.�`TŃCD:�!�|��(��o3K�W�>\}+���K�G��+���_���B�tO�Y[���������B�Z.�p��o�yƂ�M�����WxC��"���xB�49��W�W��<	mEn�����c9=<�u
bQ�����s󌸼�v��n�%�*���E@�����̋�D���co[
pCX,��=�����=#k@'zeWT�!p�� ��܎3//�y1.��&��Yl��m�Q���oi����ʳ���߰�UN�#����bhi>���_�V�f_���Y�U�t]� e�2�9Li��9P@`�A5V�Y7��Q�����O��W��Ab >)�h{�8|^�g����Q6ч��n��f�lY�Y��IIP����d(�fe��P����W1��3/��y��o��rx���apOQF�{�D�ë̇���Do�����N62\���I����g�kS��ëv^�*3n /T[�1��%�D<IUQ�D<�9��!م�Te{�%�CĽ	`�o����hR(}�B�����&�
���0q`b�×�"��ԃ.����#
�?��/�ݨ4.��"o�B�4���^���2�:�Y�1�|խ�6�B�/�lE�˸�┲|�~D���{�Q� �(����lO�ݙZ���Ns�I���یc����*�~N"�z�=�sj\O6�"���=��l�9����T������s�w�o`aV������ �R9cD�a]��)�n��y�L"d�����&_:�8���h�N@{���Yp�f��ч�l��(�Z6��'��3�:�N���(�Zh�K���A�t�j	 �)edḽJ�X�(���16?�&j�
�n����Ҋf�<.������N]~�\�u�##�`q��61J�܈.��I:|VY�-t�!��c&R/$Ȁ�y���:�'-�<������B�XxF��$^���_,]]�?)�W�w� �e|�l�xӃ���}��	�I��Um4�U�LC����߄�H
��S��D�;�u	ݫ����@:g��[KII���� ������`	���ѭ�����_��U1F��J�0@��)狰��|�E�:e	��Df��v�����������E���]�&�e�mMCj����d]�"�.=�mᘘ ����N-1�YHԛ������vG��w��|�SE]os97���z}m����sP(��f����yU��䫲���>7�H��Y,��6K�6����V�����u\Fi韏��4h2F���C_y��gzD�k��K(R6j9@2�/�����}�A���͵�%����g��XIrb$i��{���u�;9�b�����{%�%\�"���1Z�M�ۊ���� 	��� b�XQ\�Q�/��͐�[��j�H��U_<�e*�����+++�\گ��]c��A��!:�������쏄���O����-�E�bh�.4�8�W�>��m��=���'�����c��L]}�|�_�"�<o�/�8��J5���&",�H����:�E��@A�'tP�	Ff�}����+��J O���p�[���4/q���	]7�3aq9��"T�g%��d�9�_���q��R@�چ���^t��ϸ��z���K��i"��l��q���%�8B�yYZ�C0��������B�{���Q�O����bp�(�p=�u ?�Xd b!fIf0=H"׾�aW� ����љ�=v]�PW���ʤ��� ����$}�;,��<�ʕ.���*'	�XL	�T�*���|�T2f�T;�����ڂ:f��Av�N#��s��_@[�M�m��<���*8Pox'�U�4}����O^=���Y�{��}́)�}��Q0�vƓ��4�Io9K������<�"Zm�#kV@
�?y���矼�AT<J}˭wjH5�ҙ�-����ᒬ�8��ae�ǣ�B]�ʓ��R��K��Uy|�����"D6�fsW���g��j����%�?C4V��P�&��ԥ�Q:�O}�@G��}%�K�m��b~x3�nl7���MqG��i��H"H;s�"Jͯ	я��F?�O>l.��<^~28�]���"K��y<2�t�к?\t���Gz��mY�ٚ��R����/+�s� ���n���!1�!�̋�}�5��D��}�o�4Xib�f����)��B��*�� b�$�
2<�3�_�Nt�d5u�e�����3���="��sOW-w�%ۅ�g�s�(�mn�tSw���������x�i�J99iD�����-t�~s�95��I��:\pRs��XK:�w�T��2��6lyJ�vt��K/�
���+�/�����/�|Nb�o|�'wO?d���"�C�=W_Ա�jpt�r��[7��Di�����eaP	ٴ�T�V���2�jD�??�i�LU��Ej����?�����t���Q}�We����%��@ �xcw8	����X�\dJ(J�cs�����h~,-�r���r\�~ɍB�'FK`�gK�A������T�h��`��-'X��(���\�
�n!�)��餪�V�QV0x׭����R(}u+��������o�wR�_TD$���FIw-�0����-�«��W�9p�Y����ӉZ�c� hP�����5ml��T�ת��v��p,��z��l��&djJ���]Ĥ�yMMtCCC��'�o9Ҹ#-Y�8�����3��)�k%�lm�B��n���))5� v~�Wݖ;�0Z��OʉE9}^a��䎚*|�Ӟ���z\Cq�N?�X���Ċ��y�+�Ԓ�hP1)���o}�b���h�m�<�z�Ѽ�F"���O��|�q���&:�m��#��o������]*�ݒdz�O>P��魂Vg�μ�w}�~\j��d���:v�s͕ţ��H�A�*c��?Y	HՁo1�sBx�^���c����M�x�������:�"BBA�x�,L�׭���Y�'�����r5�B�Q����8w�_}�r���́_u���z�mN̥�{D�ſȟi��$=e���I@v!��ܮ��dN&ޢ՜�fȪ'����m�\�
�Tl���nu�?�tY%p�g4��0}~����� �R��[*ܦ�\&w��7a�����e�GO�f�c�48��+�>��?0�Ls�*aـ��u�,��+ޛ6�Y�4���d��7p%���¨~�������	�zKr0M�ރ��]K��CRF)�R�
����?��4�O�o�9������o�n��n ��!�9D�+4��4�)��G#�a:�I���	�r�H"��S|=�@z=��h}cv.R�؇r�0�1��I�k������0��M��*�������������)�M��J�er#����bI�&���#�ϋS����K�b+�{Q#_ԫ��\w9|����w�0�V�d�wުW��@�j]0��7������&��oV�xk�4�u����_�I%h�_"Y��0w���~�m��b!�K��1C��+��e`�3���E����|�	��5��EP�B�ʷ�b�`v�������H"�H2�p�p!>�S���~��z[��X�©ߊ7حd�W]Be���u�7�T#�Xs��X#��
i�Vc%��a�\�X�Vթp������?���Tx־�P�?i� 9��9�'�����/�
����ޥa)�G!,ϒmF�P?���$�,]@�y�+�eQ󡽽/0����-�<�l~��g���57�q�s���={hm�}�`}Iz�q��#4"�K�������T��0��u����/ة�}~&�V��N9qs\��oq~��~D�X�.Ǯ���A�kĒ�*������&�V�;�:#�cTr4���܍���ɧp{/����e�УR�Z��h\����7k|0�ü�A�H+k�z���S��ܦjbX�S�KK�����X}\���|.�T?=M����N��o a��@�7�&''Yi�}O=6�Qf#]>�t0V|,��+�y��>�������18!?��Nӵ���d��n���ɮ����2�Gy1��۝�d�t�m��}���s0+���v�/A��}B�mx��JZV��Jr��$i�W�9�u�,��K\��$�L4���bD�Q�,}�Y���E��;��¬l���Ȓ�I����NLFc2���c~g�B��ɿuuu�0�l�{����_L��͆x;~T.��NON��lc	n�*<����\��v��{�G�[��<Wko�����w�`������Eد<l.:��GjO��J����o5q!�m��;~V�;��/�ޤM��G8��#qv�3�<,KE�ȰC&����?Yu|?D�'#R�����Wq#�c!�� ��f��T�a0�W�0�$�)vf9�:ڕQ��6�� p�+���@�&7�5?O���H#Z��WGe��|���؅�lC�n^__ch3��1b�/�.!PEO�\�l�ͷ5��E+o��tf·�"6��P��|��5���3��}�:Z�>uͱ?�|s�:���|���E���)fg�<��W_�z�L���	��'�,�	Z�sף��.�`߻�#"ʈ��!���0�~.m�9�ß!y�c�^m����~Չ�xO�=Q�Z銨���r:瘍�
`4�ߥ�x��1z�����H�xT�l�V��w�k���ZO!akgf�A_է.՛\��'e�B�9^8��b�l:���U����M]�Bm�p��*����^�
e)�o�ȹo&�~
Wj�g�K�h��[�z����aP��Q�@m_��"͜��I�fi��w��	z��t\ ��#q�y��)��+"�x�V|*@�;��~	>�iY%�[%����ͩ�7�NՏ�k�3��hk�;U�5�%�5dv����N�b�737'���`U�wed�m�>��e�m��rs���ZT�'�v��n����Z�%�M���u����c���u��&�z�,�:6�.a��8�nاD�JL-e�uև���/¹+����̷�r��h�غ���C�j	=�Nt��]�ga�ں�v\�Y���.�骎C�GՂ��3q-����G%lI��S�
Y�4�ۧ;�&%�Ƣ\5�I�.���<З\�ڣ� D���ZO��� FD�iN#�"_5͘_�$u���(����0���\T�G�lX�+�p�/Ow�Yņ��s\��"��|�G�/���Y�"x*����j�>|���Ŏ�@�Ȃq��I� �W�o@�������+�~w�� �i�7�%7�A������"�]ވfM��\�>�3�Ưg����ZIz�J{�Rأ��g|�4�UQ!���Vz�2n0�)WT���������P����/�ƃN"�D*I�!���DX�����m%��eX��Z��� ͻ�ܓ%s�%�u��d�u����|��!��aј5�jF���}�E��H�U��^5���i��UY������%%�L����P������'�x��8�� Ɖ��ts���1}�'T�E���Y|���͌\#��I]ގS ����g����E��-�� [u��ۈVl ��}7NN��1|�'���,�}I4L$j�J�����>mM���ʋ�����B'�T�ah����`�$���_���^o4#/�g׀#�~�A"�n�~,1�2r}"`m��fŒ:|�
Zb9�>_85�+S(���#\��0퍝`�pVT��%�w��
��)H�H�w���ZT����Z�Ԣ�]���sV��yGϠ�������"cX�%�SEf<��ۈ�M���ܟ1���|}�]�B��Ƿ��>��}HKf�@�cNW�o����E�������#�ǆe�΄�*�b���^δ�% a费��:
=ܿ Vd�����(��h��H�qY��nYW�� ���L6��P�I���9q@~bs-!xm���*�e�Ͳ���~z�����7%�ۛ���o?�6��=�o5��2�0���O�>�|�� 2�b��1u���W��w�m~����LC�?���Q)+��r��|���\�f v�$����������>��֍9�6�v2#�?�sv�-�l�ڭ����`�7���|Id3I������z�kGߗ��]��7����G���Y��K8�#ސ� �@Q��y�	S#{p�O^>�!$��r��\<�I �U�������Q� ��T��1�r�̀���f��,,*)�	D��۷yVU^������C�
�� ���������ڹ���2}�c�����V��	y�W��k�&��4���j'�x��ဤ�r�m��">�; �-t.h���c�#G����; �*���Wb��ϊ*�c��?��#��G�u,/`>-H�1O:
�(�9��(E4,~e%�h��z���X��B��l���%�#,��+�Jņ�f���8�� ��ԩVV5��
ִ�V��p���_�2�\Q�ٸ��Q�=�򱺥z+ ����f:�)p�����|�eTUa6Lw�$�i�n�C$�Cww
�ҍ�HHw�R���Cá}��y�o����u����{f�k�����e��u��y�(��<��d�X��Np�[�E��T�d	����?��{����dƮR�q��S�\`@4�|m_��ל����=��6�S�'ϰ<S
-��h�<:2-�%�>��Yu��?Q�������qw�i���q��_ՙ�S1�j�e^���%Ӻѷ�D��9M.�P����}��ul��FX�\�����GGO�V��,̟|�HS�ϡ*�Z�2tL�<��'�}���_�����5T$��E����'��[n���i_�o��9�h��<�k�6�3<��6U�%5O<¨[V��s &�<�`/\
�i�b��� `��J�߆�K��$X����y�fo��7ƿ/���n6Zs4�3�6b���Z�Y�+6�Ǵ\�C겋���umC��0Ye
�镯9t���я�tg���k���|:��]]��JA�t�LYbf��n�����W�㓓h^y_�����BqN7�*7�0ާ7V�X���V��T0{:����a���	�D����dm�wc��%�7�U��їgU�	�
��p^�~<%b��7Kx�x��_'���{��U�)�X3M./��x]��ml��W~�՞�[e'<焾��e�dB|�|�����*1 &x<%$�]	)���|ݴ�AZN���t��)����?Z 5�����묢��8��0�DfX�!���kV	��SQN���A<3��"8��5L5�-1�|�b�^Hw�,e��3�l�c �q9'RNx'�
u���X����{Eϰ�J�a�h����.�ϔc��EVJ?uCGiIJܘ2���3Ѷs�ul���M���%����\�=B~U�� ��@V��B�wM� �P|ن�����&hy??�� e,Ff�.�u�<W�ܦ/OR:bY���xqY��3|�o���5��b��d��'��M�rmP�d��>M&@-Ԑ�I�G�|w����~p�YKpӄO,|g5��TA"A��y|y�!L���k�f<�.�͗y���gz�w�����n����.K
�j�n�9�kf�7r�Q$����C�O��φ<�(�3C!f0�헺L�2��R��}ۓ�o>�0˜d��֗H,�� ,��?!PYE5$�3������js�6�ߔ0v��~<��Ҵ/��r������i�1DU��T�Ř�#�zBB�F�o��gRBn������ƽJ�Ӛ>�'9��Fq�'�ѴC�˼���ׅ*�>�!����O�+2&Î'��<�ܤ(>{���r�V��,�q��"�>��Ņ��`[�D��7!���ϓ֬�F��/)�����l?��g�}N��v�K���]eP]��GP�q�~ܶ�I���M�X�c�6�Rŏ�(����Ē�����)q'�Ii��X��ؓh	��D��W���~�F{w���W2?䙂vĻ���z�Z�������V0�!��C��*�u���J����za3��}�����N\��&'�����*|6)��<i�V�2�"�bA�&�?8�� �BW���~lm�+�\6��o2��V���1�<����/�o~繯��|�+��,����R��g���h�	L�\7����8�s�?o7���|��� �+�`��JZ����.�Cm>��/���kI>�n�߳�7�������Dp4�/�^h٠�� .Aclhjv*u�K0N(A?�5��2�u����Ӝ��J�zfJ�vhZ���f�iZ��nyC}z�����^��Pf-�w����1���m��b0j�K��������t���v��{ގe��w�	7��4Ьȼ
߆�OOs����	���n���M5�@�=?3Y�ӭ�&������kc 8<r��*�(:����Bvp��*�
7��혉�4����ަ!oX�is�Q�\�ا���n� t.��Ǟ.����z2�u�V{�Q���X�i����M��=�����,GD����d��PB�f��s'/��v�crjj��l�P{��������w�U����2��NF�1��Y)L_t?�69[ȕ;�`aDQ��:��G�^�����S��U�ݣ�*��P��dY��G>9��}�����>X/O�����͛����Tv� =�7�}o$]廃���W�B��w7��Y��> �|�n ��f�{
���v���������8aݞ������z=��0���b[�\�W}�1��b��L���_�߳k����QҐ��n����sb���X� Ot�^59����#]�T���߮�k'�|.[�uF���]u|����Ng�����Q�̕�},Ƥ��>&�������e�#�>�E�3*�^�-.|����/��6h�������OK�_���K�':�8���p�nڨ����Q�z�(�h)����!g�$+1ƷL�o�5�rot/ ��'[-�S���2Ja��y�<���XW�V���^�x��҇��q$�d� �=j4�|��-��|h=����c�����kjhl;d����CS��g"��D�_�/G�4=���j/�X0�(G^r��]5<l��~I�#�P�ipEiL�����'Q����/
2LM�����%_��C��OG�4����+��B����TM����P����_�p�a��!5�>�N�W�⿖��4@�.�󫈛j����Sm��?N�GQ._~�kyĲ�����p9Sd��N��?�U>]g��	E�(��dJ6$,��ǫ���/�m	#*Ar2����r%^����B���Ɍ>U�>)�Nr��� p�L�N�{��lrɖ*�����2 @
��d�F�qu����'{(���Y{ZW[�rL zr���b��t����:�D�"����t/л ,s`�6�#&�+=
φ��D�'ïuy){��0}��, ��WP��@��?wn9y�?�#8���/4� $M���{�/歎���eH����?�)��7x�޽�o���g�	O���z���+��S���䁐q
D݇wE�0x��NBp�!E�Y�O�c�N}:�E1�g�$��m�1͸5�
ޤ�Y���7.��Wl��&����W���D����������z�5	�c�m��1g�c}zi~>�~��t���ѕ/��{���Vo�D�K+����',z}�v?o��,bwdќ�N�Y=x4ǮI�le�4�5�~�����C��֏���11����;�s~����"��|n��J�� ed%�Sâ$/yO9n=y~ZF�X\I�齗k+�4-2!W$�´�A�V�G*~5�,cY��ݙ���{�*ġX�~�+�����G��3D\�P3�����/�$_'��#"8��q��� �i��ܰ� �1</@�VMc��~T��g��jy����'���g;Pa���Y��%�Z >30<��i5�����!kK���MUt�<�
�]������9�h��}
נW�8��qҖＫr�:�#5�Xb����pV�U?5i�ʔ,��e��c�y?�����}�ȉz�רZ�'�2ؒ��?S�
�BZ��w��q�߮�-U�(F�+aӶ�E��5&�����|��l~�M�Ǫ�vz�<ն���&��3>��
"��������D��p�a,v����iA|999p=_�/�B�,��- Ɏz����k����O\�ݧ��(����&�t�C5�A��%9fb\ae�d�������-�R���r���ѥ<:O�V�u��N�z"��}�	�*��bλQ:�.�����`ko����u> �s��u[�[�׏l��wg�MM�x��O{���YV���ވ��SfYw�P.�
�v�w�)њ-�ּ�z� �X9f"�:� Gc6��N�T��Z�-S��b_֠Aj;v��h�?�bH�B)D�`f�u�p���M���PT�D:DM1�7>(�z@��kX9�76�wjD?o������ԧkP�HxJZ�zݫ�%|w��g(S��O������x�}
4��#,|��@�`F��h�YW6"����Q:_�ji�!�ó54��l��;[�e5�j]<...��#S<<<�}�"9b�.f�]�#D�������1����(�O���OY������ƯS��7麸�u�6��#������S��)���F���Q�Ϟ��U����&�L;�̼u�/:^㼱y���jX7 ��,�X}�m�}����$�;��jm�X�s�8�����ln��'nSv^V@����vӧ��l��;Z�B+%���R��z���rX��C�����7��%���,��x�>Z�Y����A�bWۗ���2j]������k��rzw'�޸������x�\=�d˧F�3�s[t�tg�q���9n�,q����D��:�����M�l�_W�#�:��<��ӴD霹P��`2�u||iyYE�n�sI��Q2����H�+���:�nc{P��~RB0�w�<2=;?��?�U@'��s�m ��'ͦ���XQB �MTj�y���<;�s=��k���Ч��sP���v��%/���)�.ki��-��>��r��WZx��
Q0N�����=��J���zF��hԞ�|��ۭ����^@�6����O��a.��Ŭ��c1���{0;u�e�,���5����$���	��䋋�T;��n�]&-�*	�L�����ځ-�j\Ѫu�*�� @^��_�:��P�����I�xv�>Z���Ug2�l�f����/��Vu2�[8)�ql5����8XX��s?֤Bcj9կ�6s߆e��|�_��;������[�BH�Ȅ���!���e;�~��O&ޚ�;Y��c�����/?��퀯���{���Ѹ"����t@@�¿l�~ߙ�����i�P�ceXJ��$>K� �,~v�T������\�Nt5�m,�0��f���q"z,��X�K��J�y@���`��!�J����Aw���6��tt��,�j�Ƈ�ŋ�r�[i���zE�EnRw��P�D��=�����!_I�d"��T���""�<#��WBN��=Q�eN��X���YX̴7�}�@�*li��FQ�#��7Z�o���#��W�-�u,�S����D
�<�g�no��`�.�2�5���{R�T�V�~��9 �Pf��3B�L�}zz��qjq��p�>auJ�=����w8^�6�!�+8o���K��(Q��ag}R��hk���c�`Ϟ`�^�� ��Q>$0�*�>���:1AQ�W�q}}�x2�/>6��������8yT��୭���,<||��Ck2zUY�[��<U,F�q	�導��Ƴ��lܰ�.���RX��Y��<��`y*�RV���%��}"�D�׺�|��R�b���qcXl�-���k�w�bqryMMT@�;�,4�9QX��D��/��}��t�@m���˼O��s���&TP.oL)�a�C�;��h,�~�6�Fu
���&�.�/�O)�����؍��$�D_��cK�`���4S+0��y��Uf��Q���h�l���$�҅rĽ��uR�w���|B���lu�;�^.{@�p;�:E�?���i��V�ߌx�U�1������I��1�j�!�)�]�3���YP���#I�j��eNV��7�#�h��Ԏ�|���5��h�t����$�(a�u��Ky����`_SK�ʊMTL��r������p��r��lи,�_����F����YX|��87UU��Xk�gՌ����Ja�f��|���סMKy�������aT<�V�T�L�̞2ΏB�?���[���{�%�w��S`"*7��Y<��J� ��ayy����6y��/�)�ttt������:M�A/H}��G�T�����aU�x�*!C��X����
~-��pՄ�V�20d+�@O�Q\�M���C=�A��D�&�H(�&r Q�˽C�|��NH��7Yx�I�F�D��k�v��ז4���IDŭP}ʲ7x���`w7;��K��S��H"��|x#���N����$p[�o������b]�"N[Q?���Ґa�z����"���Taʜ!H.�[~�6Z��P�c�>5��m��E�Vu�5r�8����C���9o�����t�p���,���Z�>|�Lk���T+N������ؾ{SW � W�Sq��7�`[���6��r����N#n�ԱAඬ�`��.V��ÚĮ��>��g ڃ2~��f�U��lB�iM~�(<~`�#���<Ԡ��+A�C�
�2~�st���f,r�a�=gDi||m�f�;(Ң;F�f�=�~�K�9|5ۼ�Fb��Q�(������3K*�X��&���[�%˟g���U��#�-Ǜ���.w�R[�W�H座&��===��n����Z���Q���;t|��Xi�9��/�䲍�h���~���w���>%e�:8�ޤ��"a���S�
�u��5���WGK{gUXD��%��/�=z�M	i9Vҙ���P	ƻ�\A�搰n�k�>3k�rhXߤ���������;�V�*	F�����<���iI�䪢"�Uf�[OmV�1��k+%��Ye8��ȅ,������g�T�Uϝ��\�ŕ���f�:-(�s��(y�jN|������O�UΛ�b�4E�RE��em���0�VnK��ػ�s��=��S�ӛp'A���Qt�㭨��jِĘ�����;��_F�j,���C��{���;����N��^���^��
|�w��x���V0b��A=Ekձ%c�L�b��`�%318�����@m����i�B�%{�ZZ'ڠ�����̟��6o�����UNN�%s�J�[Z2��.-UӚǡx�P,�.�}��_��S��wA�pX6N䠡 ��$�V�;����q#f�%��n}C����.��ض��u���g���w��bi�jo3 �c����I��("�/@��s������6�^ŭ��8�"/eo�g6>Aa�7 ��ir ۃJ@� �d��_2J^_��]\h��v5���9}�	�{+D8y0��v��+k��YO�8@׾�ӾJ4	�u�&�I1~{����-��s ��y�U��C��\��@�T�J����3Ȏ����^��yE���L ��lP;�8���{�i��18��Ih��\�_y����DC��`c�7��<�����[��@G�򖊜2= vZ�N{�4���E#>�O�#�va	�ܜ��]�Ki�=+c�/����w���ވ��G�'�7[��
�{C���t�/��E\@>Ń&{yw/��j|�W�xL���ϴ�e���ǨY�P[;����Q�Lu8��A�C��/�Z�E��y.�,]��ea����Y�2n���Z��хU��/�Cn+���'��8e��m�A��3�F����IB����y�6�x3`� �;8SHw#���Y��Ǌ��� ��ʢ��<b$�At��2�K�!� ��D��OȥNt aNP?_~��qj;���d���Ťn�V�ex�A�Ņm��S�����j�s[��橚�� � ��n��=Vs�ws��Ǚ���$Z�K\^�[w����R�K5w����˼;a�vc�3zS�8�룺r�wZ]Q�A	�	���Os�L����U�q5�3i�h5��Ldx����G�ֺN.5���+�����ݠ  Z�Ƕ�ܷ@��SaS��ٸ���O_5��x�@�(s̻z������43�Z9J���+y�u�rBڻv>�/8�VDx�Iz僜�i0�r4��l_�c��0���WTV6�u}�H�R̪�wĿ���9<�����W����,�`$��'RI���1}p[h�UǙD�lg52U�JdMud98�t�	}�DQť�����ag�6Y'�+���P��d=��\��&����w�jp�=8��ź*?`���:v������t~go3=������=#��4>�mI-g��ӓ������>"·Ԇb�X>]��z�O[ ��!�M�f�"�����'��KX�I��u%U�'?=������V�t����d�
��ހ�a�~�����(���\`��l����IC
m./��ס��3>>��}�~����x�?5�.��S��8߉��8D�J�]�[��0"����/j�P�֟�돊����W���Z�TXi��Hs�w´�N�_����;u	�	��LLL�������
a�AT�/??�*���B��
�w������_D)2[��]Bf��>h3�ե�r�Ԣ�E����V���um�Qψ�vS��U]��i�KC�y&�5�� qͫ��" '�q{��@��o?+�Y	����8����#�'٦�ǲ�4�ػ����^/����.����3l|1��@�!�~����n޲�� R$�f���?c�}R��5�;�Yis�8e�݄M--� X�ˠ����6�>6��5�P�?r���S�<����d��p���N��H�U�Wc+[{b�2��߯�(M�^�Ri:��3KL��R^4�H͒���(�~�9B�aI(p�����wz�!w����4������ [!s��m�_$5M��Ѭ � }��QIĞ(|����g� ��|�p3yp��w������Ҭ�,#�E�dZo3A�ë'��e�֭�������lX姹d*�b�/�ܧ%ˁ=z�����;"I,b���*�����P�{�!��8��b���@���ǲ��w-��6%']�b�(#b�=�V���C0�����w�o6~kѭl��O���k����v��WVj����bU��Ѓ���q&� M�Ծq,,e���.�'��$+��6��CT\�¤�V��l�
m����Րq~[��6%�X~�I���d�/�hx�"�Z�t��{�y�2I����@Mw��J6A��'�����j��Z��p�)��)"��KF�[���;R$���X���ς��*U �&2���8�{��C�ZZ2RY��/߼���9=}lf2�)�r��tn���=G?�^�G������א�8K�2}�Zf��ld���X����"�2������S��wD��ˇ���T��k8�3�����cV�(����y{<p��s8Kj'E�p�e��G���7ԒW�TQ������<!b;���Ō�˩w8J���xv�g�Ծ}���?_L��;��Z��8I�;�bxz�ȥ���I	��	�(���k�)>^X
��6?������蜌jS�Z@��U��@3�!iN8$*��o��-+��\{�p�c�V���y��ț�6c�w�qO�^M��%���r� 1D�J��&3���^��i%<�:~,���"�.M�>�A䲬�|
�>~ȏh���7и3��jҼ�Q��|ںrm�!X�Tӹ�[qY���!�߽�� ��n!m�� ��ht>�'%�F�L������	�����:F������WxŪ*�N�+��D�e��VNn��WD?��M��ʪ��J,�W8v�=��ܓ�2��u��]��>`���6"F�&��l�=�xd�A3.���˚Q\$xd�
F��8x�__���}%L���H����Y�2�f�tq��J��GO(�/��L�$/'��ʞ��z{��v���z2=��wY0��)m�)�P�X����D
��.��?+�b$��~��������p���������K�ȭ��b��#�kh��[w3Z~��-i�-��V��{G&�4C�۱J���j{�*�NE��j_��2�t�V�XT����_���|n4��۞ڼ���Ӆ�w���@
T%e�@8��]��*(�Z��e�yYM��)`��I�r�8����Z��JX%�9���DGl�y짬��[������ʹ}���H-�m����ɷis��{܋�}�U%���}d@e�9��۱��XZ1��2�;���0�og�ķ2E"F��Ix}-�T����F���޳`3�B�֓WM�(�~������m�5}'����_�߱wO0qʓa5�	�nps��枞ׯ^�yq	{�X�|~	�U���J�h��V�f[���sa���w��y����]/���Oe���P3^(n�Ɍ��/�6�`�u����&X��g���)	���`�'�!����v��IMg�$����	�5����O-l�R��U��1��f>�Q�w������V��f���`)���`�&�����v�#�q
����Y1��,z}W�I�.�m�Ky���?l���*2 V�֣Lx#s���@��~5�v�W)DFG�GH��H�_y��L��ޟ�kq�=��p��[[Г��>Z	>�;<`��d��"e��|V,�y�B!Xې!�Q���>l�}ơ����,�l�uܟW��2��� �"��E&ZSb�/�o��V�9}%�Q���S�����Lq�����t�@��1/L�:D,� eߵ��|���YZ��f���|�_��9�����;7���zn�~5jN�0_'�b
5K����i����T{�0b�o��v��@�*TB�,�1��2:��=��hɯ_�x��5��(I��zg	�?�ZS��l�4�j��Z�ɗ��[����d�1�8)f���7��?�R�r>��=ف��3)���������\��W��`���Ad������w��/��w]�/:���għݼu�B{��w6c��Hr���>�*����}��$s�ٗ"��{ϣ�4��@��lFF(�k�Y�D��u�s�\v��fZBl�Sm�wpA=Ϸ���l�g�hOо!��Q������)�����I���*H�������D�i��]�!�хO心��F��p
i�� a�D�W,B����P����2��Q���R��Q�~d~{�e�R�Я�'�ML1���-��z����؝4E�D���(T@J�<v��<f��#��{�kr�mK�e���&��%�4�w�%�"���	�F��M"r�T�gxʸ�?|ѣ�3���Z9���a��.�b�U\��������~J.� 9*g�y��q6��K����U��2��&�G���9biho�����?%���!^Aˇ����^����lu�4�YO`�����O��
x��������ۮ�:󛗟�2�ajR9�ͳ���%�
��SL�������Ir��k"Yc��\���`6~����κ�U	�,4�ʆ�c���s����d_���M��|�����X��/�J���բD�y�7���۸ﴩ���أ�Lux��������x�2��l�j{^������(<��R�@M{�a�QR�/z����l~�|�6�����>D�	Nb@JO��r�ui����S��Ə�P������<�&��oL0���I0}���>{�U���K��31�_@�3ʓ�v��-I�%�#6+���&�U��j���a��/��\�*���J����m��\t��T&��㏱pL�vrc;�Y;���#�c�2Sm���o ض�K�����a���"v`=�=p�7���� 8+~~�z=��V�А�a63P�yM�sq(��ny�Z�����=;i��[�?�����Q���h3����q���Y���y��$l�֔��_��L�.�D��M� 15�ڽ���bd�ǿI(�^�#�����\u�e]9xr�0j�3��LG�Qb^�
ݤ�dt�ʞ=(������&O@�==�߳�`e��?u�mߛ��~�iCL�}A݆!��҂�Q��	*$êߵ_LX��4��6r���Ծj�����H��o
�խ��6! �*#� �N�5%WM ��	�
���_w�/ہ���f.'G��|ZBhj���������P��x����{�ygۤY��{�G��he��Pr�^�	AKK�q/�*x��I��^++㶟f���H�;�Z��f笭���_���Q6�����3D�'�8�KR��X�4ʛy�CNi�wEE	�(�x��>ʅW�����t� ]q�]�JR�ۺ�"��qk���-���f�<�dg�j���?����4˗�R�n�?UA}{W�p����(��o�����?��F|+`DRs~�o�X���;=��k��+�?M|a�DGVf$^�\�`�=��0,�%l wQ��b���Qr��-[h,�!�����������-I9@~�­<'��\��xț��ar������"��G`[�W~)GzFF�� �/��qO�^L���_bk��&�
�������H�Fx_��]�i��9	��}ۯ9�c�c�pK��@={�8��K����~��v��qƼ�ֺ�Ož���-|Q�a��~qʭ�6������df~�A��^��mR�rQOՙs���'��x�<�!�f��ID��<]ӯ����tB��nq��Ч88��i���S��$ �2SR(Q�6s�p��u� ���Đ���S����yp;hI��ܩ!��X�U\p�ξb��og����c��l����1�J�8���W�Y�@�Λ������/ځ�Y�b���VdBz��h�,�HX
�B�/����QY��+�=��t�K��tUܟ��&^i�ݣ�j�.{�T��b7�	�}����O���N-,v�z^��u���u6���:z�ôs�����A&�ǆw�%�YIqV��=.0���(�� g��|�����a��foCO
=X2C�5ɚ�2�YP����(�Vh�/��$���!�!G+�1@(C���9oX�n��:ID)Iæ���X�D=�m|\�����s0�2|Z�� w���J�p�a����� �(:..._�k���̓�j�]e���W��Nt�t�p�P��?�����Bi�S^�0�Fr�d�y<p���a���Zn�X�*,J�����ʕ�T��?�O���y��1��+Iw�j�ņ���?��>�եd����WUou|�ۓ?��p����)�!�l��1N��o�\��)1�m�M=�±���ò�4�����Gp�\�@a
�i-��|���PxӨ�c˴x�O���-�-�7�^=5%~.���	/�QW�M}���	i	�����ZD�缆
-e%�C�m2C�ƺ���6]
�<_�J��ň��oU��@�b ����ye�G#/����mP���E:bø��L��S�x�1�e��is2A�s�U���C�@	j�vɺ�xu ��1T�E�E�5�����$����$(5A�؅����������������p5M����,ȏ۪^8��h:q�:Y��&� ����b*�{��Sw��xCju�xC� 8�N�=����SO��������1p�S���,��G��6~J��V�k>m���&9���ZTbF�2�2�V%miQ䖼����Z	}�x4i-�����I���8W�3�&���U��z$Qh�7�����TY��n�Q�"��<��Yl�A��G��M�l��_m
o~� ��&������<�4�����	U[]�G�_$g|E\���EܚF����*6c#%�)o~��f��a���l�7Aԋ҆������r������̗�@�=�Ç>qj�+I���M1YK���W#ÉG��
��m�&k,�9n�9����5��v��X��"R^hԷ�v|y)���:�>+�R����A��=��������y���z���J�y.�����0Q~$�s�����>L�F/`�!���l�E2���ѺJ�JEӌ�Cǩe�����D��$8:�����͘]Kz0~�)��Ŭ��?�����u=��CW2�ه��G7���Gϰ6�/�o>��]��j��%��j5��F�M����]�.��$�u֠��c�����K����j�7�2#'٢���LIK?��g���.��@�ՒZ���c�5�G�HV�J't��ilF4i��� �5�����S^B'�D��/Bìv����'� ,���m&��m�C7�9mgy�X �S�Qh�p|���v���쬫G-���X5Ҝ�5G���$��2���D�l����}���)$�Ȳ�Y�\;�(�p:��(�I�zx�;d���<N>ȋ�j\}�_<}�z����kQl�8e{eu���!��5�$�׻E�9A�D�����j�^λ$��O-�t�܅<x��˜y�~���R��[\c#��abܧ���+42���J��/$��f��<P4�e���\�8ON?j��S�3*����5׳���z�˲�kNpCQCC�Wlu�@�/Er�U�p�l�lAf��SEd�o��f�q}<����H&ِ�Y�6��~i����mg����	-:_w})I���dH1i|].>'��h�L~<�x�J��� ��UBv�.���z�1J��q��]t4N��q����v��'�q�ol<�Ȕ�@�v����^s�<Ӫ�KM��-��2@t���[8/n���H`鄑8j%�З����(��]��P̖d��ِ$1��U3[M�"���<�R�"Dr��}��I�u��]:���\1��%���1���sP�Z���� -ʘ�Hw_̼�tZ��|�Wj57� ������ ��M5%�BP��s�M+��&΀�)����V�S���=��a�R�{`i)�ŝ��-:^O'�u��?�[WGfhh�4(�ؘ�4�ǣ1��{�e��W�Ѵ�&c�Ke�i�D��'���Wa?��_�(`9IczȾ�V��1)�L\�B!���*snQ��>h��a�]cJRkE�Pي�D?�˦�ٙ�VQ��>=L��7�W[���9���!6Wz���'�Z�wM(�j�7s�MٕRY0��6|:9p�Y|��O%?n���Jg���i>��<���zB/Y��J%�,�缁;r�9�y%[=;��~���῍:��5���I�|����A@��p�����AnP�<�R5(���͓�G��.\S�y�H�f@�����L9I��8;94�$��ˁ�Vz|y��r������v�	��=�L?�cυ� �Fi˨���^x34j^@�o��!�G�j�	E��Ȣ,��*VV�N��z���q9'�(DL*��v'X�CJ�T��G��SW���Ō���U���+6Y����[7K��>���k�iT� S��t{9\�����^�r��r�0"Q�!����ͧ�$l.��3�E��k���	/t�2��"���a���d�`z����mL��(�{gW��~�l$����>Zխs�U,���(�5MQ��g��wy�q�E)������F��Mt��U��|����I\پE
�	L����N�zB�{��n������C�c�M.;����/S;;<p��1)|6<��%:py48F961�FL�~]8j3��փqW˪`�|NTggKv�T�2^=�8=����������Z���i%$�c���G��v=�zihq	;�k� hs��ݚWE�S��5����\?>v�q�҆�����J�*��(�"��������C��3u���|���!�/)�5�q	��[��VJwf�s1�1�,��d~��Y
پI`��2�_M�Z7���!7m��V;��%�F�m/�G�0{����L[��@���{��;ѕ�3��̵+7����vA'8��'ײ��>����4�� }V�RC"gjH%~��[c!�nX�xρ���q��B�3�n����̺�ϐ
��;�n�i�1�E\�����I�ͧ֑��@l��^��	����L�I��88�[V��l�r�]�BZ�.�*C�h��gK�6Yn��,:���O��=���l��\<F5�)�=�g� s�����3:8}6O=���N��?&՗�����*,Ϳ�lӪ&��I�Ƽ!��|ꑒ�W���I�*J94OS���.d�R�5m��{Lo�;�h��X�,#)M*i�i��F�頛A�F������Xl},ON��l⭁��Ėo�z�a,0�1��/m\�����<]��6i���.���}��d��.F�&팸:�\���*	J<�-��7��D}�R���$)�A6�FM���u%����Ew��.��+��eO�:�&�V�OjQ���=O~���9n�Y1A�x�R��/2�l���ُJ�Fڝ���$Ɲ�;��;�g���A!���q.
E=�A\Ҕ��(�mp������٘�m嚻���4�_ȥf�/F�jx+�����\�졿�nа�����6���C�#�<���v�ZX��ɯ���U���l����D#�g����i`I[f^ףl�=%�Ɍ2a�_k%�ӫc��ݬ�mY܅'=����߼T)ר�0���9�yg�����%/9����%d��*���7�no��/jrVA}4������V�e;lHu�����1L%z���$��E%ߝ,5�bU��[�T ����c�~%���-c�c=Q"��8):��ğ?u3��AA�f���⦿Y��9��Z�Nt��5�|��8/��
CJJJ�'�7$Ǯ��E?��ywV0�e1I;+�I	��V�^����{�5<���Qy���a�=�Fd/��o��Vv���|�1��xo𔺯P��Q���L����y+D]^��-��^��S���V��k�:̅��ւ���l�`{k�h"�T��@> @�UP�XW����G{:���#�3WG�Y���{p8O��K��?�+�W�R5̻��;�X��-�X��_���Z�i*���ݝ����jqn%���	('.��M��2���FC��FÐ�u.���rt9��ye"W�:p�
�UP��~w��Ck����VB
_Ϧ߅�
?�B�m�eQ�0R4���r�,_���@2��S����}G5\לM�1>F����6����X��6ʁ��V�w'�M���z_�n���i7������n���Sb�����n�Ut�jX��1F;���b�����|��n��]�s���&�)U��piƬ�����YB����k~�����<υ"�L�����ԇc:�}#-�d6ߴ����fv�h���ܹ�Ff�P�HǑy�v=��S���h[��3uR*-�����i�J��5r�J�}D'�	���d/u/�j����(��v���3dد�ã��˓�[�*u'^���2,���A@J����	����$��n��e���A������������.x�㬵�>k��z~��yI	��C�iD�RY$�bu��ܜ/"�/����Z��e�o�қ�lM>l^i�,�ޫI>�ն�+�ǭ�����������6�j��o<=?����\���dp^��쑖Ο��]]�0���T�z"D���|pP�����5�^��{w㔜�6�@��8_T��
�����=<��p�f/����u��;�U�Cv�l��\3:cxؘ&�B�;��͑��������na9ws�qG���J��bٛ�e��n�0/�(�dqG��H�`iǐK�n�����p��Y�I�L�XV�2�}�0x�Nm<�.rx�O;G��;�j�!"!�k+�~݂�0��xU"Y�E3�kx��81���ȃɹ,"
m톶B�1���C��s]�j�|,dh([��<�:�7QV�CQ�k��+g�$O'�.*jy�]�1�t�1	�_x��߇p��y5�[�Հ{G��z���|7�oC���!�4����C�H,�a�kļ�V��3[*��J��~��3a&�����7s3��
w���җf[�!��YL��kD����ܛW����i)�!0�r��is\pMNE���gjP�ýV�7�}�U�|�]��j��&�m�˰`��u�X�ڱ�G>Rz+�Fc'8ϊ�:s+ۛ<�8p�9A��ڛ(���Af��畾CeY�zw� 0F^�4|�N�{�y�T*qlr�%{�V�q)�:�(=����yzg�F�G��kJ�P��K�>�v�4Xd��e`}6X�Ou�7��g���7�VĄ�����&=�7�����K����<!�'5�a��¤���o ,]�����C���3s#���7�{i*���� b���[b���o���hW��PZ��_G\#&�̺��_�/���mh�6�k�}�	�7g���`x!Т2�Hj��!��൤��m��+^O ��E��$�y@@@���F��y�ݟ�rQ>�hiko��Nԉ"��<�����R������0[�;0t:�����ygR�,��W)J�rka�?�lq���+��������T��"9����o���xB��j�sG����ׇWs��U�4���HJ&��E���:�E����w3�#�c�YK-d9j1�S|��[g�J�w�֏�t��!S&�.H{5�'(�"�r=��D���!��4po���͇�=�]�q��13�aA\��.�;�����>�'�e�k뙧�� ��uE['���7
B�X�"Ja�3�1b�pfWB�p��p����Aw��rS�k"�˽�$��r��;^�Bu�2��h��f�D��ui��~��C�B�YI�i��@
# /Evx��Z߰WlӪ��=X&|���d |4���9�$U���W�Zi�����I��y|� ����pv��,�0h8�n�.��n<d)ȿ�����yJ@J�)Db��lw����o{˪tX�8\|��C������4A\c�����Dm%H�Û��%�y�*�<ǌ�<*`�K&�~��y���L���Q���j�����|*iG�<��H��E"%8�����C���	�	��G[y�V��C�����,P����4�O#~C^�(�7��h�q���Z���a�I�)�(������c����ɼ�ɨ��-�W��pW����ڊ�_g��2r���|�� �*[�����7f�c��Y2��e����If�c���T�-�;
ƛf{2���/��2�-���yuY<,�Y՘�1B�3,��y+`�	�e������;/�xx�N3ws���h��B�,i��c�\�;;�&! ᇱ{�GS����[�j|u�Gǚk�};�ܦ�<O�
�F���=vRh�)��M��ᱚX�kҟc��PжR�CKn�2θ/�Q@#}n��23�[�G���A��68��b��L_����Ӫ��d-5�A�2�	�Tϵ߿��ՖK>V~LđQJ����<9�*{�^��|_]UQQ�%�� �0���Y��'{)������Op:�����<�����ú��y±��)�W;��Î_#Tn�:Z��t�
Uh�I��"+������j��$LZ���\j��� ����	��?Ə�9�kMn_�P�+k�^<�r,M�]�_@PoB��qR�DA�b<�`*Lb&|?00�<H�^?H����k���h�:\9�k�e�����z����p���M�Q�����v�ͥ����Oz�K�ٺ��m�׆o� c�$�AdS'��qӰ�&��X:,�o�A�IfM�F�-������%�,�S�!�`����0T�T�Y��D(���'�!��S��ي�)y+�gA��ݖ����hH!�ċ����Ra��h����$P�?C~���Z	DX)w" %��N�*��H<3n�A��11nƑ��k9��[P0��$Μ����#I�]vHcӳ��a�����X���E���<����9 K�U��I���r!ޔH��n�4�+S@��7^?�q� �6L����3��p��ǌ�q��aG���F=a�r߲��2]ei�ql�1s�	����v�>��"���s#� � �,�YYs���������dU"�Wo[���WRq�L%$n�6��xt2��$%#no�`N�yq�!<�Z&z�6A,���jc���
�%��+crAf��V'�͢^j<�e=��_���P�Ǵ�B:���d���?��o"1�/q��q��ҹb��kJ���{$V��ͫ(z����'O�J�M�[��*'4Ī�� ��� Q�BlT�i�5���Ս4C���+��a�>�k�"���S�P��ZւQ�j���Q��y{"�����w	�B���n������SOS�(SJXE?��iy3r3���3�a8���?NQ(�ԝ(�YW���������"x㹡�Y��G;[�F�y�~$Q�4�5[<��^����'�������ٽ��S���x�S�����K}���X�����܁�N�;\��:��a�#����<-M��,�E�^���^��Z0T�����= ��ZZ�����֘rYE�cȨ����&������@4����������;� �p]���oL�6�8�q4�414"��\y�<6k��yjzm���Jy�~6��C[��B��~�8����ʸ���{�:o$�1~��k���®�D2�����!jV)��Z;�KNX��Vȼ��x+��V�)���� ���,� >���뵄�����(!�� |��u���%��?����^��¸�6��P �ڋ)4Ԭ������)zªG>JL�SR{\{V�2+�~,)9�65��{��W �lEUU��"Τ�椮wt���H���Ep�cZ����z���f�o�+�O�9�\+�ΎEI}�>O�'�e*�ij��Q�P��Km�� KZf'5�ہ�'���π�/z]-�4R`	m��뛟e�b>�'��a��|$�u{�X/m��,A>�z>���f�<ޟ|���{;tN� 	����Jf�ۤ��UV�,�窫���<� �NkV��I �5�E��,Ņ����x*YR�2`vG�����me��k���0��~ٛ����-�S�f7K:5o��[�:��>8���p#K��\���~k�L��\w�1��
�����4��$�|q��D�S��2���m�o�TaNE%k��]�eҀc+�o/*�]#sSѣ��tF�WO��<�&��b�>�av}���<��R��E�T����q4b�;<P�ԉY���97K]p�e�o�_s-T�c	�}��%��b��8����,j����z\�?<�?�����y ���sv�"�b���;�8���;5Z���a�w*�f0���"#/��8
�A�'�
	�{���4
�������-:��I���d�(��M�]�ɦ]h�Q��-S8~u�(���ʓ��Y[����Z�L�"o���I��w���ʾ.`ބ_c�>Q���L6��!�c�B��+��3Ǳe�d��w�4��Z�Z?'�3[�Ωab�j�zQ˄��d����>�gK�43ߥ�~n����d��OLrk�(��ȫ��I��ׇ�?�"������y��x	�;��۵tXt���f���$<�D$|��s(�f����v�roez���)z���Sv^�败�ʗpv��=���+�%��ǭ�h�KLu��c������� Gw���YB��|*
��N�ҍ������q˻�S�M��n�dٜ;0�P���;�:o��9��<��*�Zy�:<��?�1����H�Y����mM'w�����2R�D{�u#����\������B��n�w)�zY�/bu�3_�Uy79'�{ﶪ���Rc���������[Φ8rb�$���'W�~����P��q.*R�����c�ڳ�G����Z��2h#Y�����=��T+�Õ(=a��kzrA#	\�@!�z�[|�^�60��~��a�f�"hL��R��o�����>VTT(f�	�J�m�B��yr�/�\w���i���G c��nC׈���ν�M���B{��X��ޯM}j\2S����ٿ��_�kcd�:��g��ml���S����T���qS*G�v*Q�j���]�q��uY�;u A? �O6kDA�j��ﾉ�d���q�A7�<�ڜ�Ja�����V�i�Y�Z�:�]��+�S:��Ӊ5U��S�B��q[l�Ta~���B�S��_�n����|��5cK����j ���f/  �5���3ı��;W��ؘF攽��_������YX�d��"�˸.g^��n����ŋ�{����{F����xi|�Ъ��m79ظbXo��V#W�����1^�=x�ΰ�N���O?uu�C �2&-��1�i�c�c��Ăoo7����!UUU�Qr~-�_)9����s|�"zᣅ�
f~g1&r\D��_��ߥ�w���GC�'02�iǽ�^��K�ra��Ҏ7+q"W}�m*�@D_DF`_�S �si�J��R%���Ɖ}�,��e��u�n^�G/�åN��d7Oם	r4�tq�}�j�M��­�0��-�I�����7lQ5�u���D��lGD��2�p_�0r�Kԯ�+��f�Q�e9�v�-œ	m�6��B�����/��q����ty�\d�Qo���D�r���s�$��ڔ��@���6	~������Oh�Wh4�(��0С��}'31L�깋�����[3�,ֽ׷�O��Sb��
�m-��B���O�||����g�2tL0b&j������f:ݲ�۲�o������o�"G?
ƅ_T� �_^!�P�h���S���>������ήO�Ϩܡ!.\�2|�+��(�����46�k�⦻���l�vG�VF��0ț��gu1�^��0%BR��W<ؿ6�ݢ!��OM��L���J�)΀�.V���������A�'�� 9� ʇu��!��\Z�Z�'N�.�$p�遧��Mmq��}��U��"��i�֜_2�6�ܓ�x�,���C��?���U���������V��Y�2�K<��NM ?���.\g���7��R�Q��v��h��呭���Z$ֿ����un��[W���@��T�q�|���-��=k)�C*�|���")�G��Y���9�3n��z�$x���D�o�\�]e��fQ\L�g.�}���(�������k6A��R�ǝ� ��ϭ�$���hVu�&��V�#�	��A=yh��`�C�/а�����o&��-�!��b2�Ȱd�x�.!hJ���o�ı~���nL�hg����sQ���O�k)�j���>\�b�lki
+K�٫~L/��2T���=��Ǘ2����ug�Х��6-q�� go^��A��@/����q�9�2_���f�Ӳ�� �ji��u��v3�=���J���Np�����-c6�K3�_t����R��-�c�����7FU���Eh��K:��G4זS,F����DE:�a�3a�#74��}�b&qR�N82�š ����?D�wR�&g��-;;C���p�e�h�2vgg�V�"l�>Ss���s�S�r�y�K� ��:B�����R�ps�Z������!��_ݽQmQ*����u�����Qoc�J�e"�(k�d%���r�����Z[[3x�������r4쮞��D��S���I<[�e�d�1���������SD1l�LΌ}�
�|c�d��˗��Zz����	?�r�<׸�/o^��c�r�F���f@`�Bg�$*�[>#e{�,��"��U��Q�#�5��"�5Z@˓ �`�k㘽%�NБą�cS��N��[��4��|����>X\{7�D;%��8W4?������/���B@�psC�A}��7�������"�N����_I"x�yP�>��!1�������ڻ}JN�؟�ڐo:S#�u<�ӈ�h�ϵvv;�L}�Bծ�66B���k�4P$~�E+zM����9�2�f���pX�CW���V���q�����gX�����NEnw����90^��1�2P-�x����Q�8H��ژ):������bǉ��;sw�^"a��ʨ�Xm���-ʳ~� �GB���.���d/�)|��I��w�}h�gr�g�KF��;��=��t�v��ţ4�W����DI�B��,jN��B��Y��Lmv���kd�=�W��T<C"���/���@�# -�y8���1su���t7R�8�+�����{W������,�,��H'�:ﷻ��w.\��m%�a�T����g��n��1{�f�{I��v�7�^���}^�z|*& �t$����hko�;����bἎ�����Z^�c�,������f�'��� �*�7,�d��)�!��$�@b�j�hp��L{�#Xkldw3���$�..^W�C��L��e�S4�h���	�����{�>4�gS|�SN�M�{W�ۯ�[z,�[��8M�a���>���2�si��F��.v���T�5����$V�k��a�G�=[���͍��B���V����V!G�W�؛��e�a|�!�X6!l�����}�"���!�hgWU�M��L�-:��F���>�0���t�2��~ReEA��|��C�w������:��!+�qރ]6Q���Jn-:�2:�1��xa����5xm�R�R���_�/ϕ����St��W.��G���֭r�_�quD��u���`)/�A�����ۘa)�I���������i<��q���
��e>i��rvs]�P񥺷L���(�:����3��B.�������T��ܒ�	������0�����`�~�˼�S4dG�5�!��f�b�{��ƈi�r�?B�ܳ��6_����4�{r��;,.r�sw�I�K=OѦCb��E$(�&�GT�Æ+n!�dF%'�ߋ6�L�<���gӬ�ޟPUR����򰯷^�G��I��1�<���a�X��>$g����rww�o'����SV��½nlM�~I��_�5*&��9m'�{��C��|~#I4V�'P|�J�G�'Bū*�&'��͞�ݱ�,����%��G--�Uv��PL�~B���a%�&�� �,A �h�EԷ���h_g�MKT�ط�:������`)����Q��l�b�k��HdT�+1@|��~��"��c�}(�S5�����ڷ��>�n�\�7�� �HI�G��{���ú�SJ�'u���gJ�.а�����VZs�Ke�)�/�S�x�_�s�ׯ�~��c�pcL�ٺ�\�:���!��%�ʋQ�@ޯ(+�����V�<�����V���f#����귡Ǹ�l�nlX�l��lᴗ�Ƿ��BB�����{"X_��X�T/'����Q��DW) �O@��H�4�^�0`�h 
�^Gou�P�6�߾�@�9f�[ў��(Híp�&���xt2�b�>Nrņ�`�������m�k+"`h:�g��{����)^��w���w:
^B��?�0�M��K��0M���r����z#�)���ڢ
�z����c7@*a(�� ��K�A!Jȴ��x�W��w��M�}�ABѻKP�C�r�������*�{���5Ӂ�J������ی���"V��;?6^^.�$��;vgz��X�/I ƣ� ����Ԑ�f��q7|�|jRy.P��}[�{/r���(�p�];�ܓ6$�	q"gK3,<T�0����7�;0m�u��_�
�ȇ/",����N�l0�0:k����;q\Ee;��1cotɩ�L'���[��.I�8o��j�݀���#��� �h��i��@-���y�>K�}g�D}��Yʟ>\LZ��"��/�;T��ϊ.ERC��&r�M�-Z����O\���uAc�c��:�U�fNО �jɔ�W�P�~7��������++� {��gS�ѥ��s'S�hX7q�s�ѷc6D߲��(�뭇��A�Q`*�Ok^����.�����!O��2b����<�)��U��X��#����|��|��e�@k�C���ڏW�C��X�/���ΎM����`f'BB{{�Gg��]at��qk�.؉}��~pX��q�s��B�] M&��Zo��;B�[0�Z�\;�nDo�#���E4��T�Z!� zS5� (W����ݽ1�{s�
p������_���yQ���;�1Ҫ�fqM��3|��+y��c�fs������NMc&;On��_	B>��sc7�T�VJ/�5����zD��f[yw/I�����9dd}S]/1^�t��8������g��6?�1���8�b�?�2�Fp�l�V�$*JI?��SW>�@ݶ1^��~O���q~c�Px ��ʲR&HT�GN����vbS�8~�^��qBH�qr3Il�B(��"���޲��u�w#���mO�E�P��� �å)P ����׃�?VgR/�j����d��`�/����Fr.cC�3�d�V��~��}���/�8��=P��g�qQ��k`f���<�Fw�1@.������m���  �<��'y;#��k��.�L�����U̵�UضC�t�v�_/�j�XTG+�c���^4���ͮ8-��o�� ��ST�y7(i��̇r!�R ;A@�E$���w��W[)��^����9�f��Þc�,,~�߬G)�>h�yO����A���-+��D	ģC9�l�9��!���/�V�I�vq⦩��$ߥ_�ŕ�fT�-�R֔iJJ���M-lP�@�AF�M/IU�[/����ҡ����M4x�\U�x:_�&c��6�+	���VX-��<�厅A�����ֳm|&L}4h���0����ȿ�7@����.�~�0z��ɸ�-��}�#��S�k!D���U�A�G�^��$D{_���W���<Xm�=d_����YsYQHdx����v�&�<���1mX3�=r�'ԍ�������@��@�=,O�����`��l��&[��7��\�����+�����M��X��k������W#���ND�{��O��P����7&DO���p9�������M�"���$Cy�o�m�Rubw*�f����O�Rn����z�nY�-���&w9�A�3�r��_�<�gf��Ty�"�=n!�N�Q=��d�:2�����5[��9I���Z�&����h� į6�s�M�:`!v��� ��{Yr|v�#'�pq}�E
7��3�z��tE���^x	�L2�~�,���k��Z3Q�(�����->�,[�0���,��Ib�׭jq��yvb�,��
�rkX�r�x#���z���e�jKɉ��l>)Qd$��~�]�rp�	dd}�s4d#�Oe��`)A�@'��t��B%K��d��������,N���e����%��ϴ�O3(�~��Bm��ײ[������ʏ���5Y�x�J��=�9<��sk�h�9�)Sx5�7{�C�9�]�ő 'NS��O.�g�/Ц~F��i�2��%���Upv^C� ;���a�k�
��6C[����}���od^|=��m)_-G�[���ԍ��Y��� �7~Y�vNտ�mՀ��X���cW����
�L���Y����FR1���b��b�q+C�?k>�$q�������4��si�E'��g�t�q�:*��8/��vYEMU_ki]a19��6�JW�b0:���b��w�S����;�!٪�9�ا�$C��Y��1P��L
�� �fd�VI��7^!�t`pc���!�jf*������WjOS�7��|7���ķu��2�� }����qMg% 9���4BZ�
������+~SD������k51D�4��W���&Uo�Z�K�;U��4�^_�C��=%I�]���9��5�OO �N�X�A����y�y�[�=�B��E�'�|5���J����O�u
uN��l]\��Y�p�܆�~)�W���C����;g�?�d����Ӥ��o�1�����qۏM��ͣ!�mϵ?ݢ�c�e���յ
HT"��*�B���Q���FJ-�ӵ1�N��#��� fc�?�(�9��ΐ��2Z� �,αςxˍ���2̽E�|�0 ��D��`�1j�Z�y���Į���=O`�seU��ҫ�:`�O�^SZP� ��Ce~�W쵹��`���M�����M���\o	^�'u��#M��p��ó�%�?��W���3^�SL��~���Ϋza$�d��zv�ʪ�X��^g�*/��$� kv�#s��"{����Jѻ���I�Wº1�3�d����x�U�w��*.|��Bճ�����	��e�7"��G��q��wK��b^�y�g�1^9r3r�?����QϿ7���N���R��Ԕh(2w�\+�Μ�l>�OI��a�wY�?U�;�R4ZΝw����ү�;����^w~��j����ZS!5�;�k���Ǣ���&.�6�P6�+�
|���:ZY�w��&��zج����MT�mrn��Y����?7M����E�M�/��~K"~X��8�"mx������k*g��~�~+�����^*m�#��,�pc3x�抓?��\��(KC:2L�\�"ٗ�&	�x��_��'�5�͈�_�ըB�㊘l�W�wg�BܰI(����Z���t�;��I��~�W.�Jb r`���JQ��H��^#�����A�ǻ����%\�'ܾ�,��b�6U.��uD�ǝ�g,!�G:ӓ�/���.��se/11Zǃ�1Tw�F~uPy:��H��9�;m�{#�����w��cc���(�je9�����Ɋ(�~{bh��1�3,1�(�N��d�JV�#伎;��i��@�
��M��c�`9���8�ٌ�*�.m�}���I��*��P�~��q2gex����l���������C�\�!��x� Xp�� E�Sp����q�����Z9���&�hW�_7�.&.���`揁��&�/%,^|��"���Ûw8��!�Dԭ�Ж��Ϣ �f��:��w��/�Y�
0��>�%���@�F�W��|w0Sto��bd����U�Qb�������N���F{B�����4D�6�"�੶�ٓ�"�W�Z�m���b�޸�v挿��w�����E9@�n��9�͔�A[8
r��&��fdl��I�Z��Z�5�Z��jj��*{�ε��am�^��H<*�Ύ[-NT�F}]U#;���2� C����(�]�z�@�W�[��MPT$�9��1��
s��1�i����?���w�� �J^��Օ��9��۔�:����%�2���C��F�d~=����QF�FE'- ҉�2��&nw3(�����P,Ρ'��Z�v��%���/�F:!3�B���]^���l� -�002H)
�Fs�IՁ7�6���AA��ͥt�M&�z��g�L¶$�����σ��Y�m�I��%?�t�ߕ�זFG���'����Z1s�
Q׈s��Ÿz�n��+"�W�E*�uSN�1���S�>���X���gѬ2���_��=Y��τe"�W�����G�p�Y��]�����I)Nr�:S�(g'�7����I��v����)���y��E����nN�pZ��?�D)���kخ��p4:���TZ�'!�3)^s
���z�(��H�$;������4ڊ;mȁaͥDR3��a�\����yU�=4�	�_�;��I���EUb�����ԏ������#��p3�0ȹ��0��������O#-֠��`	V_Ԅ@Ehv =6�:�f��p�9W�ܑә���o�s���G"��ɨ[�_V�^�3���q�^ܜ���ZZ�RWzzB:o=���o��3��=��s�6r&[��	_J���vu%�_�!���x)3��,����Ah��J܊�L�)-��+�p���'�}i�:� ~��0Qd0u��<SK�_�Z��SA�[.������[�"y/K�����̷ii#�vӐ�e"V��U�!j�b�)���2]��~��=K�tE�����U_Nܗ����o ��_L"�jUkV�)����P�D1����=�_�	��$��Rm���<X[[���ʔ��9��'\�z���S����z|+CU�S�o~iS3��ia�O�p��V^��B��x]�(����)��ʏP���z�q��[���+�}D5#�v������Y�T;�K0��-'�2�l+��̻!P%)�oDP�{B��҂i���ɗ�"?Z*I����ň�u����E��:�-�@��C	�H�:�,���D�1��s%�y�l0�|��o��<�%����9w�y�B��I{z����J�o�[�<hg���"|Cq��Zr�f��~ZQ��� $�nĮ�� �m�������[$�MEQ�^��6?�}�o�I�aW�۰<T�`Q�ݭ����M�L��p�2����ͬ�	-ނ[7UQ�v�-��\nߔ;�5�W��a��`a�8�PL0���y���ֳb�5"3���(=崋uc��`qL�*�	Οͺl�p�Q�6*�́�lqq9)��JE�y���ZX�0
 =�xB�:$�ĝ�xyy8㰙/..�/&D��Ue��nS�{��O�Ue�/m
ѾW��ͳv0\�\d��?�4A&�^�k�9l���g��I�y�3φ�����CT,,,%�U�ԕ�n�>JV0�ݳ�n���e:�Eʽ�=���0X�_�f}��g�yߖ{9ݎ<v�]<�����Ł6�0ʌ��7v�W��Ύ
�㙆�+���F�@ddwǦ������tj����%�!ؗ����e�,�ɓ�W+�{��lx���ht/��J��~8�	�_�ۜ��60���{�2?n>q�7�w�wR>��D���?}�|D`�?o:�=����{A���9�t�յ�h����"�;9�%D4ז����Yu�?S|\2Y�Ũ]��y�ͻ�*1ۂ&)9������[��h��]��|9hf߱v�Mf�8�[����l�Լ2G��S�P���NEe�j���׀KVl�x�`i�#O�@ET�;-���L�f��֛2���3����l�B���v�m�_�	����y�'��o��}��P���&�Awy����qj~���M��������m�{�����׳G|{.|+Z��j�4��ןx��>\�Fx��A,:�#���>e��v"��n�FvW�ju)*��K��& ���`��S�k���zy���$Ņ��ԕ���ӱ��k��=!�h--~2x2�Z5'h����V�kgGO�|�M �t���X�d�,��Tu�����9+N�����c���,�����h��g�2�i�`	sc-�N}���\��=xk-bo��BY����*�M۵�j�uN �]y���o�В��L�����-�i�]U�/�`.�}K��gR�\�Yk���7_�����k�Zy2�X���04��.`o1��ϭ��.�.V�t㵌W�hQ���8\S,QA�*n�3�.�)���b�+`��Y`��A���~�ҫ�G���Q��ˋH�ڧ��Nf��\pw�v�őd]Մ&Z�Uqd�^'����t�^7��¼mg�q�������������ü�l���-<�F�/n��&�{�B�Ы����Ij[�����~F�7u�T���a�d��B����`N��4��6���'�oϴ>������A冐�~�<p���w �ͼ���,��zaŹ!#u� Pc��	:��n`�?�,��6]Q��F����^x�Z,׺Y�+�E��/��N+�;4��T��B�X�T �*���􌚨G��UDp�5f�7�|Q;s�<���a������W�$F�q��7�4�@7��" �h���*:�<wa�G���۶�k���=,؂Q�}�WL�hp������a0"���y�߭�r���7A���e:�5��$�~�����*��Z���=�K����(�g^����l����wD>�x�Y��l�6�k]��B�:��α��u�7�<�VF*63Mb���n��B�m�%i��f�BEz��	���� �ls>#X� �.q�Ր�)�ul�kʴH�s���Q�A�&H0��;���=:��m�pQ:�����^?t���޷�N<V�l^�k����EXٺ��;.�o��zYwƝ�0Ư���DK&
.{R�V0������b�ܳ�N�׻�{���b��v�G�Y�B7k����9���/���^�	��ԉ���os�����0����%��Q)�vF�/��wY�&��WlXu3�}8%a����ž,�?��uŹj�*�'lN�.�U�,zKֺ}y�ݵ�?��<(v[IjRc��a�+dY���	h]m f���m�g�^��?���-�Q�uL�yBb��޹���O/�����&#|�V��=�hb�ǡaK�g�ӎ�Cay�p�O��Mg�Zb2�n���}o��69h�����P�S�lFlk�򿾕�8ϯ�8�5W��d��-�<�U�����]t����"���yȨ�^�txx|�?�c��p���Fق���ך�Sކ`�E��:0O�����j<M�u%1)�"S_<P{7�O�\������q%�aI+��<A@�0q�ҧ��W��a1|}���C^z����uB9N2����Y�əq4Y�((�54�>�B��l��l�se8���L�x��+'RZ{�		�Fp-��|��/��?\*y|�A+̅��GQ{����"���'r{%�zX�6��#x�E�c��J.���@�[���
���}0��-7��T�Yj}-A�CNg�NX��샩�%U��X���ȣ���]�[;���x$/F�BP�?-��4������v�����5�y�C�nw�kg7�0� 8\%���	�+Q�W-B*������͙�a��G��ԛ��!���=_M�h|h���lĐ�=T��Z�ج~t��sJ��D.���S�_��:<��E��wO�����uU��0b/3���+�FN*��M@�_��|4��o�����l���2ȱ��\�}�kE��	Z_�k�{;��3ӿ2F���%���Q�C�n�/ևH�!�26�{������Sù�	a��j�w�T����Pi[q����45����i���Ј𝋑Y��2;v��moo/���s	ƖT�E*��r@\^�a��kF���b�K&������{	�o��}��ct��&�g�-��1=f����וUj����y��� ��u�	y�wp �(�/9�\R�������l��ԅ��X��B��k�Z'r�8��Ki)1��e�7��+���ѯ�>vh�����Ha��ϋ���$ߧ�ׁ�K�V���r��Uч���/(~ⴇw��Ŭ�����@0z������w��k_o;�&�<8�i�����?6H.�L�_���򪱴��e���M��?�Wr�S_f��� !K�	���㙁۲�,��,���ѢơL�'����e��Z��0��|�	�(���5�F����-��j
Paܵ����r�^�x��������=�U_�������y���M���ECx_��к�]鉼ԃD�e����o��W ���[�0��Z�I4X�b�WJ���t岱��}�%m5E	/�
��m,�� ��jֺM#tG��������&J�K����� �����ɵ!/uQU+�J�Û��l���S��O�<�I>Y�O��{�छ�<��O����=X�g�7;Sl$s��Zd)z� Ia��ݢ���=ڸreE�~x�Ǝ,��$Ҡ?R��q�}���1��=?�x��6,?
0#�h�lԸ��y��
��R=���8'i�Ǔ	�W�]��7Ҧ�Lr�t�\�|���;3.���1ki�E�F���-��O��J�*O)ahe�G�\-�,�6��51��S�Ŝ���f����9�b��D����ﲔ�~j�=���^��9i��f�~���}�a��K	`���	5!�����-�{��vU�R�*H��M#w��C�i��P�)i��ςDRqh��dm�R�7��'��rOk�����o��,��o�&���3���v�Z6�B"ǔ�F��I�/>S'�����n�a��Z�q�����|��x墅�ؙqx�叠�Rh*�NQm-&���eF���6��z0*�QO��;��[�f�����o�מ
zi|�|����1lƳ���|���[Oi<�4���v�GYd��'��'�:�xc�H���݅��*�^�iS���
��:�h���9$����wdN�Jg���Z�����Bx݃��Lm8�~c��v/<���X��O ��7nUī��\��$��*���ϲL�M���b+�Du������m6�Ҋ\v�^��s#��)�45&,��8�*T0���*N6Q�k�YM4����{T�����h
��\n��pJW=5���4��C����Q�����Pi��$Gǐ�n��nD:��F7��g|�����{;�9��9�:�h<��� ��z2ֽ�����������/��z4�� �&�۲�@�$���D���]4')�0����x�Ym7=�E�
p �.����/��^������8��WSߐQB�,ꛖF�D ������zM��b��/K���;>(W���N��-��������d>1s�R���lIŐ��.9�Zo�	)AHh���h��<�	�c4�TΤ�7�7z�����)>��z���[,�npN��O"�Q���T;l4�<�c���k|���|��Q�[)��QpDI��Gţ��%b�3�y��e@/��������;;g9:�k9�D5XƝ;D��@��5oi���
���^����:�6�r�QZ�܊����L��7 ���V�V�.�&]�{J�s�2$��ʊQ�n��8Q����ߗ��=���F���/%���Zjyw(h�p�PV� tƙ:�p-V��o�� �"t{�k՜��ly���T�n��y '�R���u��!�I��.��d@��hY;������ew��T��ڏ��
��Ga���������{4�I��׊Ȧ�}�(

hi�%�o��N�6q��ݻd��G����2��/�'�^K~�"E��LU�� _j|�X����$�<��K��߻S���6cUa;2�4�#��{~�$�Y�?B6��v�G˅���^h���!����7�&D���"�_qYK�}B�ҟ8Ű��I$Y�z3�W���~�1��4��	�$�M%���e>���8����{Kfw�LR��������ߝ_;��Sk�����'��ӳk'�1WlLQ��l��`"�O��m���RHY\Γ���ۼDZZ�9U�[�Tz��p:WO��ܸ]�<��7]N;?�����GA����x���(������H�y��Sx��nw�S�Ŏۈ�p!�C4I�(��q���Ɵ�	P��.� d�$1����B�����^j3�	��9K	Q��<�=:X��ځ����������.���֪]V�cum�ϋjG����Z-ٮ����Ӷ;�P�PiP�<S6"ȣ��(0J1Sˋ�=.Dpn�譡l�>ja���3��m2�dJnL�[h��G�yӯ0u����x�,H_�ҭ��;����x�);W^
�T:�H��~��%�~�U��.�h��Y���ɍ8�|���%_h�P0��a�Ƹ3��!�Ci��b��ۜ��.1��@�����4�]R*�o��$�H�T����p��*o�x�)��}`7�������㾵��6u����@���j\����d׏C��QZ�n�/VO�ev�t�h�b� �w�I�9����+����:�j�*�Ep@��4��N�	�7RL[�z��x���)��FQ�č�8�|�P��S,D��m��m���q��ɥ���䢞�X[���� @�mB:}��[���y���N.�/���P�����3���'v�qye�����щ%h��V00�Zu���g���_kC�̱���
��{ ��������n�����'��g]�M\[����O7J�CI�nF1;�rQ�U?��9�S�������4q�����^��B��dyy?S���G�t2�:(�	�+�[꘣�+7�FtfgHri��j��]m�[ I)��9>���aJ8�����B�b��@�
$�G*r��L�ˌJ��S����}?�0����sc퀧�ߣt� ["�L8Ե�`c� v�.�H��@6�5��m��v�}�����y&�8�d�}*S�=�7�1+7�2�p��?u�=��V������1����\���P7�RHvo�+I)��~%�|؅�M�%;M�Oqnɬ�}36g��׳�����a��+�ԫQal��a���$b �9ݻ���6�
�3bn��\��:�G}�m,�u��܏)L��bQph9����y��4�
����AR��yR�b�O�\���,���6�իv\�r�=�=y�/N��f$�z�]D۝U����D_�����sZ��E�M����0ϡFg�N�#�����ԏ�[��$��,���1���?*��U%��>���e2��7�����S>�6\n''|�c�l�A��z���w>�x�{6�s�dax#��V	� �����M?��FyQC*1 tb�Պl���h�<6Jz�im�񑟷y��%
��؍q��H֌�����Oٛ�vE)�6��"�\5 G����y�T�1�/9���J�2�!7�}���2��Ä&�qU�΀,��&IdT`�����Q9~�xXZ^'���ީJ��R�25MX,͎��1�:�c��~%�995��°���Li.�F���{���Tp|ݪXc�7�,8b�b�Ѕ�UȤ.�s5�!b0S�� Y�w�<2af���)�HPET9sP�5�7m~(o6�K�@�m�#Bû|*�RIQt�<)�|�Q�:P[�A�3C0�&~й��?�>��͵����U�%��w�f�i����-Q���<�=Be�{�_����:Z�m�*N�{F�����V�&*�/{Ѯp��)��M������ٺ~-g�����[�V�ǿ�� ��ڟ:��w���DU�ǻ�ǗY~b�.vr� ��	915[P��Ɨ۽R�Ao�I_�-�t�sQ��O�*o��������D��16ܶovVôԤ��Qy�%bN�8���y!غ[���ѽ��I�+���.9�_������qE�rA����?3�j<~�3DAe^zڳ��-|�W@�(YR��xu$Ő�"���.�z��[0!/t#lc_��F6
�2���r�~}��t��P_�ZB�r���s>��j?��c��WtD�
 �G��Y��peN��ii)�PA ��&�[�p���T�M�
�Q��^s��}`��H%�d���f|��F�:�ܩO�T�e��ٶm�N�h�.�F���v<��ll�V�k'ӭhDf�Z1P�aZtX�	���ǝX�'Ϣ�KQ�f����0Ƨ�ُX��ߩ��}�w���ƺ��!:�t	"��2�Zw�G�=~X�ܜ��j-��{wQ��Ȇ�"��תj�ܞ��|cm�9�Zz4���!��i����[AIH�Ц&2� dD�n�U�_̪�Irg&�3�H�Q�)f�=��?�L�̟��6��
���ȤDϞ �����8����Pp�N��T�椧w��d,�;B[g�s��#�5���V^�� �K]G����r������#�o�Qj�.y3�N���w�鐹z��S�� aV�R�_���b>�eG��������Ʀ�Zo��D���Z_�Hmb�k�39�[��Uv[�����

�K�&$��?ݭj�K��3z�����4sXUh��a�����-�k!J-��zQg��k1�p��`Y�ͰM|$at����XH� {g��%r�h{��FX�C����}����h�`�L���IJ���WJ�
M)��7s��̿[Z,���}�-1yg���S}��g�0 /�H�*�R�RȍH��'�ZU�9# ����X��'�b�ym�NA+�P�)���`��?�zh?���{��8�����Lwq��6�O��$n~X���|\[Ӕkn��=4�?$�\� 8iE�шY��ƄtcB��}6����%�����Xi�L�D�0�3�M�D/ϼ�F�-��f����b��.�7�\�

�N���3��&�D� �D����HBq�B/��S����3W�����+�s�}�]L����*B���Y�o���w���:E���Rk����l-B��O8H��H��Jpv�y=�&��S!��"*)��':��2����kW��	2p������c�[��m�yS��r��Iu�GO2�VC�h{K��Pip�p�t�J]ڱ����vr߼
�1{s�@�X�ԡ�����#��)�3d~s�B[9ݎb..�L&�<j�|؉0O�۫:#��Ol;Hx���(���j�_�ڪ�8��U�̃K:N����h�B�~uy0���w�nG��E�U���_����l'��(�X" �ұ ��k{�q���}�U�ᩛ��SSS��<����@i�:���μA��G��<E�ؘ/�sM"�����Tr-�i'L��?�'4��R�3�y�.���a�_y���6���&��JR�h��� gb�\����-:-���V��������r��eZ�#���0oT9��#�����ѵ[X �o�_|F9!a���|����<{��xĖ��䊹�����;@�@�LJ*��.�6Ń�)5b.o�-_�=���W�״�i�x:713e��Sѥ�X�5�s��1~�\R����5���n��E)4^o���;�c�:ZL.���r�ςikk�Ꭹ��i���V�c����trt�ˡ#����lua=�����%�"r�x��\Ѭ����u1����e-9��Cm��(侲e9�ޚ��O���4��<܎��@_�����k�#!;#ؘ�o%�^@�*��]&��KO<��8qi"'UY�zS>�d�u�la�_�����<8���׶v�x
	tM3�+(I�;sѶ�)Ô���P�@���{�]�(gYk����h�	dſ|�O�|g|I��s�����:06_'�_5Dqs�d<G������ʗtB��ۯ�Bt�̄s����.���,��͆'=$��Cj븗��b?�Ln�u�{�|�2��b�m���$���;85ϩ��'���PM��L5��I��?Ύv_K�w�m�]�7������#n}=e��p������6�"�F\���B#�"C���^��!K�SK��Pf�"�%7A��Mt��
�n���1���ƶv�=!Ƹ
��c7�W�X�yq.��M����Ìٯ}��3����i���Ѣ�z�XBؽ��|�?�������lA)��(I����vS(H�e�J�rL�y}>q7�VJ�-��1^�
G�-���V:,����
�iqs���|ԑ5��da9g)_��.#b{��4=��������{�	��6�ȅ�����D���(�3�"������223&�4�@HS�2�����Bv�M]Cչ	��Djs2�Z�s�]�Q9�j�9vFT	�<X�Ŷ�����0���c,S�A��T���72U�Oa^p'Ml:��������*�����Dp��pI�"i6�)e���@��˯���&��8�p4�^]5���xo�F���tp���\?|r���D���V�s}K����z�GP����~Ҝ�(��=��5���Z����<��/��g ���I6��h�s���כ�6ܲ�o�ݯ����qT>���C+�u%Y9���)�Q˛��=5u���E"���[P�_҄;52��F��>�:��!c <��*����hLK�>QE������;��y��W+~�
��O.<c�ݏ�wj�n-��{(����^ݷf��'c�ZBQ�T@���r{%m撥�MՓ��ذ�ھ�#��y.j�C��5�vA�b$���m~$�4K�T�>X@U��N��d��w�}n)��{��/�>���.��*%/$7y�)�{֛��#�D�r|�K���I����5݋�9�.qp� �է@�KzO�>-I�ܠ&�H����S�y�ܰ��!"@7_/�MMO���oPe-�]!0mZ��ir�6"3��X4�#/�AU�v��l�&PF�=}�9�=b��~�ϙ���LM.��ۣG��##�5�Տ�,T�� rh�)X���p�����5s���\�÷F�
;:���Q��2ܬ�열��~,� �v:g����\�>�ᠷ:��V/�O�p��"�yil�X�Y��Di�~�\�j6���&�R�Oyi������m!v�]�*;���0�Kq� P���[n��EV�Sc��b�ge��V�`1�r�	љ^V$K���#��f?�7`p�cI}��[:S(�%���1G!�D��%����j�����綧��Oq�H���1��m��~����Rh��d���p�{��Q�7��7��n�c�o�wdJ��Rmh�w3^�:�:���jF����)����P޶-7��P٣0��#踀���z�$���P��-f����\O�G0�#��JYA����]h���f�S7�Hi|���Y�>\�p�-N�����b�ddأ�d����2�A��:��/��vM^	>�Rj�b��Ge�e��u;m_���;�`�*�@�[<��3%�]Y)4N.����uz�#����ww=�XRKl~��6�q};��k���.��y�[���ΑG�=�7z}�=	�E��;w�CXd�r ]$����W�T���E˺3��}}�Ȇ$��n��Zͫ5Z����t��,�=#��sMaX�>drZ��~E��jp*j��
�Зu~6h�߷�[;�%&!y���QB�-�ɫ'8P����M�ҝe&U��MR[:���
�b�5����*QbO.`I~{�t�bY:�na�ǘ{�]}���J�U{��M�- 1R2����G��_�jA?���X��U��t`Wbh�v�S@��҃է�����nՒ'oH���nv�}w� &���g'r`��x��z�eN��}~�^�\?<Oq� �#���bgM�AAv��6s���I���]�'x�������R��!�(�W�*�"]�	S��8�~K�%��5y�GAMT��s�(f���͎�ܦ):���9�{���~�׮���[�G0s��G[%G[%�����់l��,�iYqW�+�p�#�g�1%��y�`�P$P�d�s�ģ�Wn��4-$��^�	4bE�>\b>�U��/�Mhhg[A:�o��0���hWz[�����*��9w�]���]������VÆ�Rj;Se���(�Lz��?���҉d�/8��(�&�j`�~`΋+����rnG�u���}���~衃i�>`X`��m6<��;���N��h�MmZ~�����Υ�h()O�]y3�rVo�p�C�	b�>I�z.f@=���ԩ���t2ep�*̐7ò�K��h�R+�\��[�ݝ���%��b�Ä�y������=����~�ط�����.!�C|���r\�x���zp�72`6���/~I6rJ�������&�i}����)��:�C�Qs�W��[I+�7�`�_1��A�?رJrn��.�{Zr���<����Hc�D���׻7�cUĝ	ɳ��͍�*0����w�U����rm=o�8���?���~s��,����}�;�W�6�s-�'�.A��!l��m�s�y�ؗ�L�7�l�\I�ѝ,w�kF�`o��mh��Ѷ5,R�x�D�wi���m�Z�=b�#6�v��j ����{k���$e���k��kV������B��ŁNL<��+$���D����1qWK3�V�,�L8�߅(��m�(�/`�IZ�P�ƙ����̒��I����8��v}Ӂ-�*��
8�9�٪�{"����nU�w�2ЍC<4GD�(���J�i��j��<J��o��ٙ5�@��.c4�_���v,x�~�����ۙ��R�����鹺�	�����	�tAH�P<I�u c!Z���D"�LYQhH����I��@+RZ2V��z���J�����蝚�ob�-w�T��8O�y���|��=a���͹��?��d?� �М�<({��F�_`��u���#��(�V��g-%�z������j�y�-�;
2Z�p�M������a^Ͼ���T:�3�����r;_���':�U��"iW�+N�ΉA��lƚƨ	�z� @M��Q����81h���_�ܣ
��y�Ϋ��1�`�>�� %q�Ƙ�����p���d�a˭�K��Ki�7ۣ�&=�5�jƒ�d	��wzS�����	�?Yv����z�E�f���0G�[x�H3���}���q�+��Zq�	U�*C���f<�{S�3�au�&�l&�⇒`/'�@�:���q�A���|�K	�H�D=4J���^PT�Y`��D�O���{}���of�Aj��*ڇb�ڹ<��������Gҝ��U�:��@�>������FLە���V�d����8��GKf6�5���<F5� eBN��;{rW s���4x&~/F�)b*N|���M���p� ?g�o�F���糮�J1ny��ȕ
�K�h4J��n}Hm��:��2���S^ac�!�{q�B��#��,;so�'Q� ���5B����`��/���������6��|#���2�՜
�;o
���|�[��xF���К��A:?�EI�������)�q��ũ���$W�~Ŭ���̐R.�$�:~�p~�\שa-N�[�7���;
�U���w�pU�O�7�H*`��9��Z�a#�v��D�6,u�v�i�f��y����y�[U�yUr����y�_��?�VɆ�Θw�]l4�0#�12|ii���k�l�p�!h�)a�m�^
tB#�Z搪�1��X'M���;ݘ���0����˞P�<X�Q;4G9������ N5�h̽�q�R�;Wr��~wT²����̅��q.�f5����b7��-O�)�x_�iMn�zA}��@�Hr����r�*c�3����f��sH��`�2(w��9�������;��ђa�f��u���F��<y��O�K���)�۴JW;�D�|}c.7�M�rn{�b8��,��x����;qI�?;U�&����l�H��MUu�<�E��Z�X�'<����	��I��Z�Y'�r��KmGA��f��8�|^�N��I�0a�Vޤ������u��3�7�P�'����yX}l?���g��[��X��}�t��b�����V�~"�P�AD�V�^N/�Y�(��;�ABۀ�'N�'*�oP�N:pT�W+	���sK�q*���D���Ò��1	��Z��@����ӡ4>ʔz��/
�^���k����|C��nM��8�7����N��?sZ�5����S77�:)#uw"�*�`wڼ�gb�tF}�b৤�Ů)W�Hf�f������.oy����sH�ٕ���*��DI�bRk�@(i\��^DZ�D#r���(_s�f�8Y�:WY�y���qi��A���/��'�6�s�QM!�3�A�vP�W}�AUN��MF���ت_�pQ%�+����|M��M�7��XVU��[)<"����BK�f�G���Ό�Y��w7��y=�5�=˨�p�P��P�|OuyЁ�m������-EW����&���z��9����9HpAV����a�aDޕG��:.s����TJ�ރ��c���Ԙ����� փG����h ���xKZ�.���s�qO�Ϲ�fN]7�#��R��@�J)�s�����:�qh
��:�������\��\�O5E��S2e9:cZ�������	U#h���3Q���T��A����A]�|������#��ű�bf�n������bI _��41���}V�� �_��>v}�K}�6��;kO8{|gDnp�q���Z!E\U͞3�uU��ϙh��)��@i��% A	q/���t��U]7"�#d.%�6Sn��VL1���0D9(m�$CR��s���?��l�u,N��m�=뺈�I���E����/���W�?��|$~�\f�k~va��Q��E
��(�JT����]�&�n�3�9��(#$1��
i�eH��Ǔ�n�v�9�5l���&W��|]0)���n�N>Zo���[lzZ%�./',>$�.F�׬������ߔ�&����s]��ư��tƀ\5�9�P�DK��i�V���R��\.筎M�kX�EV���&$��~3�B~,N�I�~©/�:c�1�6�h"�I�'vU����g��o����x@��tD�*�1I�a��w��R���UE�W*�I�X>Xn��M��PW�N�i�5�<BH�����ߋ�5�6�Ct�U�b'+	e=��d��eB5�,Ӭ�BڈUR��9�}gˇ��
^��`�d��l?��}�\�1�#���Al�q`�/�N�3���Ģ��6�8y@%�@����m#g��Cc��%�����˷������`Y/JI(�Q�f>6��	��͸Uc�\B�\�~p���|x�+���������D�S�(����k
�E�s~�������ZBCS9�@�K;�`���!�Q�_ID&���$n�4�
ۑ�`Ẃ׉��+6�d�͵%��7M���S���� o$?�EC�<�u���N�v�j<o
�V!�t��O�𑆰���Q�>�y.&71)Ϥ�BU!���=.u-�D��Jo������]� ���ݫe�M�;YI����h�܀�>�lZ�;���X�6c̈���f����yxr��aD$P�z�ʊ��&n���� ��*��Kf������/kA��~��j\�D��^���{���ԌwX�I�\��rF ,�:|��!�1Rٙ����~��Ap���o#�tڲ������߰U?��'����Y^�qI�P���'�2�	`���Ғ>�J*�F��-9�2j�dU��f3=�@t֍9�Ŵ�<�y$�p��jӖ�ܵ\��^g3Y|7B���i_���xJ��h�6����^P���iw�1@�Zs�d���P�͹�G�w��{H�9ʶ����%�M1���_���?�*n�o|� ��,/v�˯��r��\�qU3i5+�5ńo�[*��V�����������-	��)N���#��Ž�n�D��.f��z�<������ϔdIm�a�܄޴O��쫤����o�4qG�Q�J�P&erV��	ei`�&z���M֟9��I��(���f��Hdu�}[�0ź���>4Z%z�l�$bg��gjs@��Y-��ר�g�B	�^o���7.pO�4����@!ta�3�MSj��1�5��j�]�V<2k��:Ǥ��j�?ЌݐK�d.#%���m̃L#:ڕ������[�Iob��{��uP"�[;:~ �%lR��mtq4v^qл�-.a�Tn���d�5e{u�6v��
���|�g�z���\�i����S������ʣ�p���vr�$+wzr��p������r��WM�Y��]~M�-!ǐl���%�?(n�}&#l&���`!D��$�W��S��L��ލ���z���#�,�
<�M{���1�*�p�׏��s���i2<�M�j.�Պ��d�.<����K�̉�nY�Y@�4�BrTת�j�y�1�`ǣ�>�s�D,ICȶ�ф�
���|؆��߈���=Oڏ�]��ZE�K��j%��(~UA:H?94��p��0�We�&�8^�q�֮��� �Q`���%�T�U�$��rt\� ��������ee��]�c��*?˷��*ꎪ�H|
5ܭ�� �oѧ�'u��-�[��N��?p��?6��/��o�~���oG
���6������>׿9�#Pߐ� �Z3��ꥮ-
�Yݟp�@��6��-�/���y���zˏB����%I¹S�Qk��9R1Pp�x('���d{p��N ���=|�[p��l)/ے��K�r�I�{�X�m�H��[��ɼ=�P�M�<�����h����4RQ�\����SE��-'����7�tl �:VCx���s�0�o4���~Q�+.�(�u�h���+��2/����eP�7zʤ���:�y�C�x�ɾ��al�[�^q$>�+�$��ƳԎb�}Wo��^�&�#,yL7�|Q��1��>'�R���&��/d-��e��ݞS���;��ށ��Լ?�K�^p��Up��ņ���AՉFآ�L��7ZU�,�������=WU�&p)ɜ�p�	�V���cH>P2m�>�^{�P��.�}�{%�M��{ji?������tUx�]� ���	��:7��!��jIT=��0,[}��>�W|:L����1�)�˽%� Jx('ח@GI½������Z$���͛ܜJ��<JY�Π/º����@��ӑ� %�����Q�G]a�B��R�C���&��"�咑F�����딮kT_���D(��=��H~FE��� �5�5�lt&K�M��j��]=��M4��$�N<v��^�)����LG4�	��]5K���m��d�~��:�;D���u�W�Qȍ� 1=��xL\'��e�j>F3��|�&�Ξ����xm���(����H�'����*��v[N�X,���7����C��T{������T2ސ���D_D�ꃁ܏��}?|�6�M±��~�X��i�Y]يԂ�=��FN�]���s��R��R}B3��^�'�eJ=��n�����2��_Q[���S8�֓�%_H�{M��o%�2tAa�F�^�rP6c��h��> ��������7f��p�-�Hxc|�/Sb̢f>�|r�����:���x�|!��cK�]R��d�_KD�)K��r���/P���zGߓs�؄��ȇ݊l� �҄���@�çU�V��&e~�*Nk�3��ӝl�(�O�A����~��7>���~k�_���&����	��GX��1��-��Ĩ��R�F���O�I7k���)�ږV)'�evt1�{zi�Q<�{!VX�P�ӥ�J��{������iF���O���!�+���V�6tRh���P�!}Jo�8pr)��=�R��Fה����F=���j��5B�t*��|k~�-��-�\=%I�T�"B��'�s��wG�C������۳�.M]�n"���W� �dC�ħ6��͇}��W��\���+�,�lH�����d�v���|"ؒ���Ʃ��n'��*!������Mc�Kzѩ�"eҜ	!Z�KT�{<R|wWf�J�����@��{P��ygCХ�R�>��#���}�lA��l���p"G�;|���W��Ŋ�Q�[W���v��)�ݯ�L)�5��v��gB��d��]y�t���P(4n�\o�8�I��W�|� �9�������p ثӕ�{(87������d�2���.+�0Kq�)�r�|\]r�M}␘vH��q�[��&�"晐�SFq�>�/U)��@W��f?�H�H����(^l���T.{�S+�8K`���b��pr^�dW�lQ;�::<U�?�^ihH�<�@���0�U���R^�bB��M��v�=*^���'���Y�7������� ӭ�6����'G������_$�s��*�v�vs#+�iHm�����a7�X+��2E��-�P�[�����g�����-��e� ����=K����:c�V��r�͔���i���"�A�,۞n�]�f��X����uhd�{�[�#k�2�zD|�4��_�h"��YD˯��9B9]�(�.r�J�{÷6Mg��+�:Yo���3=��z�N��$��2s�0B'O�9[��������%ȁ����*�覦T�̳�?9~�l&�C�0}%Y�C�_��e��<���qgn�δ�O�W�q[oV�$|�1܎��l�H�pa*1^�.}'�&f9�l�eM���
�R^4ԏ�U�.m�3��˫&a�?��Ix�*<��FX�����d�a�.Ȓ;�\�N*�+},0�JGC `{�u�2
gt�[��	��Z��+�T������[����&��@7A;���<P,P�3�ٞ��U=M2� ;V�B�	EK;���n�V��+�C�J;�Y�0� ���$w��"4��g���R����/-Mb�z*������/}Te|ޒr��pVw`"��H��@�%�Z�W����"�Zuז��aOY�:�9u�J��ih(b3��jo���E�ڽm�J
�o���e���b�d�'U�4t���:�U~D�I#�<��MjG��������A�~#-D:(�L�ԾW��ۿn�k�dy��X�j���;EQ�P��/��U�ē�6vŚ��a�^(����)�
�%��A�zm��q�)}�3bF<r��y�9*�����W�6�M��߆$.�*�k_"��"1�MeH8AcOy�BQ�FF�����|�3�bh?`�-[Ce��� ̎T؜˵��Vy��$X��;���3ᇗ�-6�Yw��2�ѓ*�����>�:��)�^	��bs��)4����<uOG8�������/���v�h2�M5��&��7�N��S)l��4�{m���ԣ���]觖3j�� ��s����/���@C�����2�(��n���BC�_[/�M����Z�J��in*% �+�'
��̪'��q{W��,�J~ji:_4zR۟�Jͽ�m�Z��X�QW��JҖ9��d/�u7��u���hj�P�D�l��Iv!$����T����E]̸��/�����2�#�^m2o�?U�q����Zn��=z.���*dODW���;hZ�&�S�H^8?ޔw�-z�$��I�._-/����	<[��'��<�c�e1 ���ͥ0+���<`��0ܖ�U9���б�Ƌ� ���CA�Ï~`��\�f��P �w�'1������ڙ'���w��|�۷���S�A�Φ��|U�e%a2]������hB�w����0����ҹ�^4�*=!��|v�8�k]V$��3��W�$��w9I�x��D�&L�Cl�T갯%e@R�+�����C���y�n�ԌO�h5�s�扶ӳB5�d%3$��8;��M��;�=�x\�+;QR���-�ܜ/˜_�a��\���d�b���%Yo��Qb�q7�Ia䨰Ƅ/N��t6*y���}%8��S�<M][[��&�<�/�Yr.���t4,��uS�>%d�~x����ji��@��������{���՛t�&�C�Ŝ#j��m��h����;�~����'�^\�ݲ&���o��-2C��2�I�Yg�hn����]D��@T�Mp1>��}��#��OĩW%���e*޹���]m�+���T&v@�^0/���]ﲬ��ut�[hN<H㇉��Сd�>�%�՛��i#�_<+ /����Y����B�n�[������}���sz=\�W:ϓy5�$�%��U8���%��Ť������U���k�(��j�ݿ��E���Z���HU�j`�����:|# =5.x��B��.��Sy����l�z��H`�#��b=��x��"DQ��#�Z��s���������8y���[<4>R>��VF0�<Q ws���M�ο��;��k�~���7M�7��T���kΫ���w<����:2�E䧼�h������p����Hź#9��`�vO��P��+�i����p?b��(�`�Em���n(Ky���\�u��ݬ����a� pD�	�՚��'���K��� �}%��r٩:s��e�9��*��9y٣C`<$����*)`n���6i��c��gc�:���_Ȏ��JP%6����[o̗��z����'Z�<(�P���Up��U-�h,�t2�[�~��!�7�Oq��M
���#�@��N�k@}��9�X���
���k�y8�AJ�ʙ՟��óю8���\�}���L]>a{l��^��n����d����Fz`/��ma9��4�?6��A�X�f�B�y�B)��WU,�E����P��6q��|�~_�f�����m�Z��A�Py$�����8˯,*}� :��Yk=J��ҍ��g�����56?׮+�P�����	�~�AȄ��@$]`	���P������-����{"��?�G�i�����Y��ʉ��>JxW[�c�#z�+R�]Ft��\�ͯj��|ZU+ːoO��'*b��}�3������5d�����+���^
�d6cTܪ�8ּ
(,`�		럯� F@Ԫ�,H��hmE���ߺ)#��a+�ǭ�\KZ急�l�����ߏ<��l�M��tՋv��ti�d�(J5��g����t��oy�2��[���^Nh�n��w�>��{�i��+�rDժj��q���j�7t��7�b��-�c�ڧ~
dWV[�_/���sa�����y�ގ� )Q{��*k��q�H�n]s��-R���-��D�x_4�����%��o�t�NS�������`o���;��U �>z,I�J*?�Y�G�W�i�zኺk����Xp�*_C�����b�����	���*��K7"7��f{F��^bI��UI� ��\��S�׍A!�ԉ�!� #GD`�5}�w�L׬ڣ�sy3��� =��o���a���,Io��[� �҉�_A�������T�#�'���z����Aav����SVlM�z��� ^yϿ5��D�V��D�I}?��K����oDu�=ءd����r$�\� 59�(߶T*J��fO��W.�
J��.t҅���У$�1��_����<n��~EC�4��FQ�W=�pzz��j̺>��nK�U!��%��Y�Ω��8�%���˚;l�\�T�>U��H
uÇ���#���É�^?~�y[Ki�WA��Pw�i����f�t C����lF�x�ߞ���h�O�՝���Uo��u�V(Rܡ���C���ŭXq�]�;w�����z��ߝ�g2������k��J�׈r�|{�"��쏞��o��/S�Ѿ�䛊��X���U����A�Po��Y���5H��2%V��3z�B$�l)�����I��;����k��j5�iS�Ǵ�.�ji�j9��▰W�o�:Yk�W:֥n�:X��H;�B�ۈEz���E��&�k5}ҕ"�H<#;��(a�����ޖ�&�D8�6G��9;|_�f�k�_��kS7@$�T k�Hv���t�`�8��w�]�:7쮁a�[����J����\m��r'O�w.�k�Ȩ�P�xՅ�ޫ�����Cwl�~�� m$x�����BHf�e�����:րi��qO����Oz����њq喾�=}���R���5r��#�8�^��e֪��S�Y`�1=��	yeeZZ�9ƹqM�4u��[0�K|�����(��[�<]�(���I�M�G���ѿS�����^�【�g����Ɗ3�Q���]��ߦ7�7��g��l�D-�-��1� t.Z',��2��Պf���/a��ǰ���N9�"4P-��3j�l�v��﷗�j�5�:дE@�Q�?4P_Rx<�>v�����BƸ��L�c�)=x4�$��H�[#����
�g�l���)� �/��{x�Ң;�-Io��q���ז{��v��f�g���1�[��	,�b�@�y����p�E�GR�uV��z|v�ldg�����w�6��P�u��Ϲ�����Zk����ǐ5i��q�=j�^/p��	i>_
���a'�ka��߮aM�?��>�+��d��R��`鮪��6g�;������Xp���|HCwU����c��Lq�ٯ�O�ܛ�6����Չ�T�Ld�YMn��Wޘ�q��r����_��%���<���"hwp��Q�(��BO�_̌}��makh���QTU�c��*T�<������&����LS�KmP<C���=..G���ݮI��L��acC��a�L��f�e�H��XoO[����Ewi����a��~�y �R^��.��b3^��u��@=���_��߆�@��3G�x�)C�d�;<�67�`�����ef[I��6_�X�8��?̖��/���v���.���i�FV�1�0���H�p#D���'xP$�e~s� Yش^���ϻ��_�:����]�1���D�+dx��]����rU3����A%}`��F�u�ju]2P�1�V�ߩX�4�@����������ҝtg�c�,+��N��A�JQ�Z�*�["���u���JUe�;�-#e��-����O����ڭ[H�I81 �,>}nEX#	D�����g��ae���o��Cr*�i�U�~`:���Ӑ1K��hRn�Ms���/�/v�8��,V_t۾"�f���Q�C5Eee�'K�q�h~��7aR�}[�E��#(SUA����5��;����I��UQ�qX1����y�I9�1����[���-~�{�!���7{G�`�1r�^��eD��Ɨf���e�}�J���ʍ�~ͬ�Y�G�o�:-���Ս��6u�lB����3��\1�*sЕ[�-*�����[����_w9��q�{V��^]�xrgC���?p/I�4�Y�����'�,Ci\S�>�%�~���+8q���F���#��#}��so��NH��9O[pD�ƭb㔛��El�(Q�ߜ��f_�)ů-̃3�UȪ916�k�\w@55�/ŪX%�/�L�a�tU.gzx��R7�dɞ',xzl�m_�I��s;���b���U|�[d[�'�6������*8i�:��%�~?�)0l��c�Kog�E5�3i���":�ٴ�d�"�m�ڄ�<ԍc���I�ros��j(6��$���z�����1wl�~��a�j��%l� j�y�m>؏�*2�'�[��~&i��h��y�@��Sӝ~�h���>�W�<�����M[(0�g5�=���6���BX��(ٷ���	�^�o�����I��6I��B϶���T�������vg���,+�,f�����U��y�`Iu��5���c	9�	�nݴ���(��q��M���x�ϙ�u����>`B� ����mUa���_-_xr&��)��eD�S��[&>
����|[��^0Ll�Kh��u�!��k���f玜���(3�q'o!F��Ʒ�'�c��_�t�UK)̙����C����|�»W(�B��u3��V >�	�8d�{	.�U�,Tj���y~��g4�~DJ��'�aȵd�E�N`*v]&ᔙ9�,��U͔g���2'��8�|C�gR׶������ LY2��v��X�N@@Pm9G�y9D�nL�+	S+�T{0.�E�~ ����2ôy=����D^'V`����.C)р���Yy�ƴ��H�T�H��-:=�nɌ�n]a/�X$B'~K��d��@N�cϪP�_���z����#�߁C,�XϷ����zneIFb�1����7�����}#��I ��i�'�*��U��!a���u��f������ij��mhZ���7��yI��dx�&."t$�H�H�� Բ�9�m�7�,�k�TL
]!��)�F:R
Y�2�9�B�/�����+�u���Aqyy_$�:t�#��_�+���ő��r�LUm������L�	��p����Svpȟ=�SH!b�GD*�[�|#���ض/����\Xx淳Cw�ϿYƃ��u߳�����W\tp�))�5�>���;m�-�W��6�zC���y�_����0����N�Vs�>c����AFH�!��9��Cy�x�������ۢ�WT׋��@�Z���h�vaF�W�?Zo�ݮ~�Yj��.��8���"7]c_�k��V�=!�>!�o@<j�9�آ�1F#���c�x�����8�f�8�ư7�GQ�G����� ��Tr��q����x/F�8t��Vy���*��k�;Nz����w�p��\bfcM�Sko�U��n�V7����J�jVv�pt�?�)ָD���n�\�o\/-���:+j�N-��J5��w)�:��L�W�-���I�,:��k�e�Qi��c�6�K`
�΅�b/g����UA���Qwy����C�d�^i��~-L�t�nX�H�T>��3~p�.�_b�mŸ@"d��п�Nwx$���5�����ǃQIP�������=�of{f���@a��RR���b��c#�\� � Qj�X�	Lt��o�LI��!�N�ZTy�]�s#�'zpQ��'����Ᏹ�[v������[�ܟ����?T��l5Z���'|��Ϯ��ȴGH<�߫W�E&&�L��ftv�i��*�F`:QC?�X��i�Iۯ���J� [jZ��y����VUw��� l�r���8�c��͆6�<�8"tы������̋�:���ҒB��쾔��1��쯟�|#~_�O�����8zGB��~u ���,��N�<oH��fk�|j�3��a{��ß|xu2�� �U��.���[�
���J�8�~�|�C?c����z],&:��_���?Egyi�շ�HS�c�QclW��y���4��Ђ�O�s�Ǐ�_�ҫ � ����`��	]�#�+�*�h��Oc�V-������ m1���5��ZӦ�<,��m`��r}t4�/<.�W��õBN���T��T�����d���:���F�蟧�'OHl1*QH����\h�Oa��U�����Bv&6���Q���q���(�2���@}���Ϩ��w�ͫ���x�끫��:��8Z��������Iw�/A鍺���,��X�L-�!J7A�t��p����1�1���E!ť��,�a�M����h�� aJcJB�Ll:u���5���Z���@̖�9�A�Z��Vq6>\�ff�v8St%]A��}X�k��78$�2�Q`*H� �n#&X�̹����O:��&���,��Qeyb(��ě��N�ھy'w��Fd�J�HOYy���_]���`O__�7�7���?�ؔcV��~'���6]$Wգ/+1#���Y���N�YII6�bΎT��������caa�����T�j�|VU���{��>��e��5�ڧ��}6�##uV 41{�0abW��������� �rE�()ޱ���1��{�����T�������v둈����@���rE�#�m��Λ�pm�qsjb�p����̡�`gb@P�DA� ���*k��E���vo�	=���Z_������"4m����Y�:&��i��|�m�%}�*�a�$�;��_1��ly����)���5Asȣ���臒�(	��e=��D��'@{@���N��m�A�O�]g2��[�T�m�`'�Ev^۶o�D�M��l<��Mf�ps+\��T�u��ؖ팊�rlD�^�;�"H�:�#ۈI�3F��)���rJ@�O+Z{D�������O;|��y������/zM(��֯�0��$(V�7}��h�ЫW̦���D���>���̪��Z7qW���H�Z�(ԁ�MN���㡡�X3K70�݇��������
�t͇���r-Dy�'FH�1��Șa;�[F
��ó�{5�xM/�"��:��a�tv��r�]�-
�#�q-#|��
��F�Β�\���*j7�=r�G�$!E��C�i��Lp�Ӡ�	h�[s�+ ���֢Lh�8Q��A���(G���Ä�G��R��,$;����3v|V{#_Y0�t;�-ꟃj�=��V������Տ�>��(��$1����!M��2r���i��MC>���\�Ș�<}R�-)�˶�P_�Z��	&�^,n���>��H7�I�p����:�j�Ս��������%�;�H
�̱GCJ�\M����1�����YQr!�߽MyY|�{��)�0���� ������C̱-'�JH��B�"׷e�v�FPL����(}�:%A�R"�_n���5T7���	�{�J�VH`��ǎ�`�.YNg�Hlo�j�)�b��5��w����@�w���S( ��kA�Ί�Ts����x��8�P��v찵l�� ����gO�I_ǈg�:(�Y �[���������`lO��<.3��76��9D�5���Y�����V=���_�|��n+v�.���Ș�~)U����g�5o�J}�"%ƻ�z%#��?Q�D�6���8 �U߇l���(��_H_�sW4��vfr �bE����2��Y�0:�=j|�R:�'sPs������nL����"�G6%�_U���@	!��3�M.-�;|?�����.�w+?I��N�*|�j:�q�0�2}W6�>�x��@vGvf~Rh��Q�����,1��`!b,[ws�R�W���w_vW4�r8��'���|��HUZ?�q��G8���������C|$"Bh�g�˓�Ƨ�eN_.�<�Ľ�%�#�t�^���]�c!fh�B��-d�~g�|�m�!� F����jϖ�"���~���Q
��[F��l��}����;��ng�ʐ��x!�6��s��(���@@�{dz�F�D�Xp8�CU�F��kd4_����9����U�ݓ���U٬�>���ɏf���k��o���%`����/�!���G�b�p�m�+#���{����!�8I��-ɤ�=�&sL2$5&*;��2�rdf9@��s
��Lo"P~W�J99�Q%�x:�s�O^��_ڳ���9|9��D����_��<�6�9D�u}�����*��	��vMpH�ϵ��J�b��m���7H��9�
���|��;eF�.��=c-�z�=�~\��a�E=��5�6p�,�ujz��X9dEl@�	֪mE�bj(ƶn��d��T��Lw?���	�j��/�A��@�[s������8|��?�K=�0��!+P�c�#�?Q���7�}�G��e|&_�\.k�ި'�Q41�tnmi�%�X�׺ :>�~g:ml�/;C��mD1M�`��O7��l����
f�^(q�2�~=��8�-3�;��d}V\П����t��Y)~ƿ;�4��~Mm����d��Ζ ������($2�w��{s��XMt���\������$pV�d��?d��0�n�+��������h~��dw�L�\j���2��6k�����J^Ȣ�g���Am����9���ȁ0C ��5�AYmA��Ω��ʎ����6�\3�� ��b���%�.���\�mG�R��)ύ ����S���j��zY�����jY�:����Wh�K�j��H�fw�í�>�3��.�¢�ĩ ��lJ�F��P(�h�cP��`R���"��(Ivh]�N�vs�D�9�6�8׽�t��e��(1�M��
-`2��*�kNSh;���(�#E��nm��`1�p�ЏͫW(�`Hv�6��:? �HT[� ��e��b��)��i[���4q��-6B��)�˖�j�+PZ^�����2C�-���̘���=�>���Ft�����k�6�`d��sb׬�Aa/�Z�2�K����oKO�\�al��f���	���2�9�8�bЄ��v�1����I�� �W^ߥL2~Mۋ��}�GgI���bI♖��-3�n����n�gffd�[[r�gH-�>.o��uR㻙Xm̆n�籓+��V�:�I\��^�Իo-S����>I}�� �N�z�|����?�QZ���ME�]Z�o>�8�T�AF8R�d_ɜ]X����Ĕ�(~#B�P�5�l�`���\B$�sx��M@���_�ְ�w�S��Yg0U!����*������3���w8	��66�a�~�y�"AH���O�kPz��#u�a��3:{��/�=��}���hQ�u�P����yQ� O�;��p�n���n�L�'oi#{�o�ĭ��`�m'���MD�
纟P �{��MKӞA��6܌�0�_�d����4�~'E��j�����?��:�%C͊��ј�1��߶�*:���N��ɀ��nͣm뙨���9�I�	��8��$8��}^��u����@��,F���M��HĬ�`Ez�D�s���W|;E���+3(�bN@ �%N/tB��L�W֍��U��}����ַP�w��0��$�c�GW��n"(��AĬ��㸰>M:��Y"'��>���Fn�"��e��>�X�?�P̓�����J�V�����Y�\A�'�˝���N��/�1
:���\Є�~�����B��sZ퇿��<_�e�i	
�WT�{I�9�>��,�l��p��yB�>6����{)L��T��$�2��q�ֱ�;'�l�;��u3��e��5<�øl?�[_���
��v!�h��ѡ�^RU��a.fT�r��L��w>/�q`��DL8v�Kx��/
���� ��|����r�߄�)΢[��4p�ɥ�{|���%)��?j��~�]��K�^ƕP;�r�5t��3[WT� ���-���b���łd�ρV`k���K�L\ǿ9� Uk�Jɘ�"����w�_�r��Z���_��"���}�����A�w_@A�n�c/^5J��5��(�(����������Cu�w8"wx=�-��ۜ�ؑ��T;B��_8��a��&�Y؈�6c��UGM�/|��M�\��<��a"ɒ TcÝ݆As���l$��]_:���)�R.&$e7�V��O�-I#�������?�9OΫy��BV_g���$O;
�k��|Ujr�)"�OY����T� �3>�v_��Jky�^w�ܯ�d���t244|��Jv(7����X�/n��ao���%�
�/=�U`�&a� ��EN���Z3�L�����V�f�I�RM_�{����ĕ2��\�g{%In<K�[�T����u�w��ԍj�ܫ��f�k�b̯��s�'d�]ɔ~��zb����9� �JI!1�5{d�Ϋ;��L�Xq6779������g<e��8�8�-��|��UX��٬�i7��w��n��j�}|�~�\��MD�n����K2�>�2��^h�/��o���U���:�� �a���ѿM����	�-{���Q�;��Sm��	�,�2570��5�t4�Z����e�$��Y%��(~Ta�U��l�Y�t-�+$���&�8����:h!���^����R��^�֝��ļ����[2�[��z-x�ˎ���3����
��ZΌ.���I�lT(���?�-�a4{� "�_:�C�Hrn����:�����cƎLgv�~�21G��(�"�Mt�ԋ�TI�ʑkK������໎R)Pga�9�?K���n1��Qb�Q����p̯e/W�r�oq�Mrd0b�:P4�6�6Y�y;mdd��u����@�⋮;�M�׋���Y�EI ����wz�� ��̂��b��759���%���+�%0E���y+;�Lb�_�h�:�'n�YԐ3����8��l�ػ��i����,M�Y��ʼu	U�[����޴ �z��˱�qw �O��$˘%1��U�=Z���KyIs\���a�AT���q�K�U����O�����4E�@�GԆ�W7Y�Z�v�~�E��ь(�t ���\-v�h������?��oOX�� 2}d$+��	&^��S�
z���W%��TI6�ݹ�Ʈ��B��]4{��ۚ�������M_�u38��Q����^�X�NJ��_ĝǪrCm�����Xꠧ}'���
�����MnN����5�@�к�S.�1�`H��*B�����q�V��PR�p��NY�"Y�����%���p�"pG�ر�"����,o�$��|vz�?/��b�����S���-Be�4�}��C�l0�^\�O�˝�|(~:�<{�8�w��E�SQWJ��i��e����#�F����e�vg8S{H�L���垹�y�o[��גn���>X��_e�m�ǉ�E��+�e8�,�w�e���D����9�N�%���M�
�Xg��tG\&�����:���S���ZwJ��`V5������`���(O	|�SV>�n�Fuj����l�t+���gt���;#O���6���I)�Q��*=L��7Yt�L���������E���y%��?�;o�9!�N����ּMvL^�S����pӪ��7&XMD�G�0��#����7�J$����}5�^O+�V��R&�b���m,��\+�����(gV�<ɗ�q�O�h~[�?2���z�/t1�)��AeX�U=��q"7v�b�L��ܱk����}6ӷ�Ӧ�dP�s�C���J�%�xv�_��i_R��Պ�x� 4��������9O�rz�?YLa��F������힧[1=(wӇ̹�[��q�Xn�_���)���gq�E��,<�����zP[x�_���(~��#u�����K���?,��������o���鵓��rp;���di�6�uߖ�,��i��'z�_G!J�&Z�&� yO�c �-��C����O�����z���@�jd`0��f�'���&ЕK��L� �M!-�
Ǻ8x��б�lW�ۦ|���$}����`8>�Vv[/������o�a�)�j��ʐk�p��ݷ���UYYu٬�mi�s�!�i
I����NŒ3m�fn8����Lj�r���?�0��=�����0G�����v`&΅�.�~���g�"�n��M�`����WY�.\�I�ę�p�� e��v���վ�/iLQ_M����d�������b��%��U��oD���(�e�1�����oL���9��f�\�FV�`�pJa8�[�R��-��������!|"K]��*''��݈�R�a��STQiN|������p.���]q5�|�¶bv�Gn}�t��������z�f^����ǰ3�.K�H�g-���M
�'*e�*I�̃�����X����Ј*�(1�7~̲�*�0��;}H4fe�z��+۞`u�������z��2�d�b���}��b�;�Y�Ԑ��������vr6��%Ec�j�ülb�vGC����Ǫ�~G����ᇫ��m�i4�H�����&D�)w���e
�!"�H�Kϲ��%p�8��A��Wv�C	GC�w;�b��r'�h���h;�DزÎb)��Oϼ���:��K��<�������;m:�,A_�I�9���J"���}!�I�i��\c�a��G�eM`׹\��F�J<�4�c�O<����`B)g���.m�T)��� U��L����R(����a=���H��"��`�}`t�`a`�)<�F�}A��b��Q�dU�̳v�e��;urXڢ��9�ja�[���i냀�f�ՊLK �T�.EH��0�_��mg��M��Os����G`[�щ�%���@�A2�y�����M	zD�Ik?3$��vK�X�+ևx�J�o�,4�M�Al�y˙>�᧛M�t��T<E�C��tV�yl�gx�/4��(�� Dc�`"o������x�]�$n��Y�'\��ci�w).�,Q������m�4����H���UZ�1�gZS�'�L\�w��H:</���� �=�_h�R��ZJ�$���e�tM�y�b���{�"���k�M�@�_�t��,�S��oרC0��J;��H*��6���A�UW�<>��Xl��U��t�_ʐ������/�&��U��x4�Jo���L�OҀLl�E8u�	]y��v��"����O��Ih!h���R������!=ɫ���.T�����=K�
����E�!p�>��aY
��V͡����1�P����4?��� i�UB�lZ��8l<Y��Qt?!�^�<1���	}/b��r���M2�m*�k���F�X����-0j+d1"�ܴ���F"�k�;,�b��'�dZ��f�V��0T�Q�MD��JA#�#�&������m�wg�ղ7�8G�z������n��� &-Pd�^$+�c���q�W����1z���ҭ�Q/��.�?�`� B�G-��:���D7�*Y���1��RJ��V����ooS���?��$���o@�F���;����˽����������"�G6�w�p��Vվ�Z���HT��¯Y��iY0�%PBŁ��J��E�Fh�Y�T��D�����9��ߺ�n�z-�J��P��`�5��*I�i�<����A ���������eN=�%I��'��n�vi��Oլ�7�/M"l,��˶�5U��cʌi �ϗ�������K��ԇnQ�oB�LD�Cc(�%���i�'��L�A
���a=A�^A�z%W	�{\b����-��)�F��튫�y�y�ؤ�3�W
_�ϐ�˧e��3����K~}{�̗��F�6�Dr)z]�ێ���>�@`�V����I��E�
����[�/��Q��Nhq>s���c@L���[��e�WM��&�K5�,��5�8:f����L�Ze��D1H�Đ�VS��.oYh���m7a"츭;����-��2ޓ�Q ���hׯEgT�O4=�){C<���a	8/�$XTm������R��{��oU*=�w�~��-|��E�p/�1�%dE�~j�}�"X����@L���Z֒��$�)�����w�hT^��.a��:޾+�|3�\}E��J{zߕbnYe�����%����u�d�zY���n7>�a��M��u9،bs��������qe_�ؗ�6ܝ{�bc�X��y���,Q��5����~�*{j��+.�y:P�R�~�����4%�Xc*c���[�?�Fݛd��g�!]"���*
�y^�yDab��?&2ꆁ@ ~���6Y��%SŔ���Zj�j먗:��^k�LX���ΌFd&��(���"ȑ�&4�N�V//wn�X�6��"����p�2җ泽t2�F��D�-�N�R`y�h��C���&��B��J��\�p�a
Г�qJ']"�@Q?#Fܞ�y!ń9�#�ȣ�ܯr�g�`"���2b�6e�N�}eK��sU��*�HC�{\[`JN~�S�[����wR�2�e�I7�&���N�ֻr4�9�|~5��pꕼ���Ld��e����e=�X>ۤ�e�D�~�ڒש�3�>u�Y�iA�x���Ț��Pņ!�f������>��+�-�<-���~�C!�3ud�zLM-E�&��&m,a&�?~���ǭ2�K���sjx�P�Ƭ4�7l_�5#ܽ��}����`�xI@�7$1N=21w'���ik8�a?:��o��)t-s�M��D�F�x��Y�9U�ґ�c�G��*�]n���f����N=܀=�ݡׯut;B��*�:|4a�r�Jv���m�z��d���}M�)A|V��%�ޏ�.dD��(�$G{��C�0�����@c�ckfCm���j�,�q�ؕ��ODW������{�xyʱ��r�t�mVC�Y[[�>�["�����e�rDI�Lx>h�f)b$�
�䄸��P�P	H�Д춵-��JC�@���H��~C�Q�K�2��Y�N�� $�����t$NC�b��i������\����s���N����!4��\����]��K�b��C���;jK�9��e�0aYz٫�/b\
2�D����ܦ�V�	T5J{�d�����"�L{J� E��&�(��m
�I��H��ؑ��_K��5_,s7/���M�*i���-M��n��p�(�F��0f�sM��^���W`	���ܵ(��!f���\̜y}��Y���������.�M���H�y��Z��r���P�3^������×�c���|�U!$��DԄ�]C�����k�Q�T ![��܃H06����5m�v�?��?��4:��{ro''CĨ���_
� !�@�!h���D�*�b=��}���:���v�?��Aod����1�*���p�t�W��6��W�B}���]�Ug�#�@�X$�n{�B����'�����k��Q��L>hkJ��Ǜ]��eљ�.���?�ޗ�ds�:���,�V��|�cǻ@�0ٖjT��&�L��ɆQ5[������ F	8�:޲��~�"Ĳ�HEnFu7��%&�I� L�@�(M:��S����W#��A�h�W�b���M�$D��sM�["[i6f{�I�ZkLo���H}��`^�Ĳ<�#�M�h�b:Ҷ�WH+c湕@�L�Dn�K�m�٥�����|(����	=A�Ġؿ��_�k���DX��`�p��9��[S1�7�Ǳ�:֛�^�.�|Tu��센v	d���~��� �|�+�_|h0ڹM\t�!��Fex"����5HO�(�~;1`��M¢�A8��L\�y�����>)���yg�3Te�Cu���nЅ����ں{n���#�Թ��q��Î��h�=�>Ky�X&�h�W����cIb�ƻ�J� ��"���`8��m�(i.0A(�@j��������vͺ/�+8�0�$���a�M���3Qڪ��a��t�/1�i];W�iVy�jS�&����E1��*�NU�2����.�����|�E��,%$�6����X�^�G@L��sU����ep>�T��+ڊ��/�O����!f�J�Q�g��c�W�UVp��s�N�ׁ�|�(}��`q�����C,^�د�<ܫy��?�t}��7W㟲~^֢���{������>�8����DLR�*�ΟTs|���,{�w�Ͷ�TZ��]��@���q���F�!��h��^/��߽��k�c�$����[GfNS%��,��_���b�Zj�т�4�$�Q�����j��>��?��}͈�lDk��)����|~���0�uob:���.�������[���K��� l:���v=��mۃlN��2Z�k�>����d�v:��c��GU�t��j��]c��	�-7B�M7����?C���pl"�yK��QkM��jO�F�G� �'1b�=�I�8A(a	��O��to����yxZ��5n�o�h�����d��)P��+���|mu?<�Q]XJ��#��b��$�V!U%1k��	�ݻ��lL�`�3?�,ME=>>B����;�#��.����U?qG���c��/��������������Z.kr�*!��$WE�X�[��ۉ���qm�oa��n��[���']�I�AYϻTй��WR_�*	Whuw[�#`;�`:��Ѹ�'p��Lu�9����;&�
�x���F݈�����J����$9��]�$����Z�A^n�il�0~��0s�G5�i�ʻ�y�ϯw�k8�F &��[��n<��M9�s���cQ��(\��0-ڣ.o�9q��(7mh��,0,�!�KաM%�0�-���$���j�Xv�܋S֪��w�z]VQw�9�ʧ�U�p��O�U<]٘WR�w�4ef�'���4Zpo���J�?,c�]�gX��{��>��}#��T��7���
�LV B��%0V��?�j3!>�D���a�k_c�eHs?v�g�O�&��7�$z)�B;��T�������~����I��k��J�Iݎn ��xa���c`F������m+�A��|%\v�d��5F+R���w<���t�"���\�{>@]Җ�!p�\ť�
#oC@��f���3p��B��L�L��d��i'�l�J����ٝ�d�X��G��H��$PMr�69��,1`���Q  ��������oO��9�p��8z$�^l�:�}*K*��{�߷��?��6��ǿ2��:�~56�D�8t��[�N�b���a�2�9@��
��H�@4V�T���7����^�W$�̢t�&�����_�
1\���1��3�xt�Q?�D�W���r���p&(FO..&��9�z)�!>��0F�}uɺ?�?�o*E_�{���1;ܫq��cG,��,���R��`�XII9���a[���-泤eL�K$)$Yl�v�&�PR���*7G��W��F%`{��whr6T��q�0��T������e�+/�~M�D�Ғ�ko�eTb(�RM�ț䟿N��F�]2WK�d��]��3`l_{E�r	y�C�;L�p�����m��FT� -!�7�"�n�_��ַ�h�E^ΨX/|������2��������Q"豞��%:
�)��S�Q9����<�~�*Z���M�	6�=��_B�����͝�ۉ�4�/�Ҭ3WR������7�@��VE��?@��ܖKq��5Y�t�:�<	��h�F�0���&��?��XG���GT~��w���Y����w�?�~z��l�_M����ۏ{�O��^lbVBt_�;a����/�B]~�HG�>�	w7`"���ϭ:��[���j׭�+���׫���紋����3�4�������<���*�,`��_j�z�6m�u�,�q����
x���P�+m��r���<���*M`:���f��D���e!]/>h\���I��/vO��Y�������BvK)؎��Y�΂�C��M�]jgf^����W+:fM.Ic����p�a�_�[��8�}��  ��j#����7� I�[�*I����L"⣣#�#fU&��^dMB���L�*>�L��L��ZX)��N��|hjĎ����E�4?�C��.TO���ȘCm�-F�0Ϋ�)��]�C�6y<g>ĠPϷ�{l�MW��㠶2��w�$�Ƥ_�+�88��V4�V#Z�2��TʢT��U꒤6��a��7�8�� ���ˉ_5�$�!:=Zv�_w�T]KΉ���_	Ձ�hj�k	X��K.z�T<���;Ey��Ϭ�귍/o�ȡV��0���^���\V�f�krg�b��t���aR�����D��ڡf�.z����@���j*d�Y�h�@1QnBvs���HO�����s�+F~�Јj`����8�L?����@Щ +����#��+�dP�x���i��B[��IB��8�{���纞"�/G�ɵo��K>�1�i���P8�N����eͷ|�T���'�Ef�f�֎��|�7A ��7�����t�$���x�"U�:�#�������~��μ����&���}Q��g��;��*���$�VVP�aݝ��xz��<w>��ﶌ��Y���,����b�jCz���+���+B�q�tNU� ��z����]Ǧ�6��`F��d;��������xٗs���}�*i��W󥹸N���Fd2�f�D�F�B(��O{w/���{�!�vb��k �[�zW8�7��?b���u=,?�D=�8�V�K��l�K��}�] 9P�PIZ�8{h�y%F����^�UcZ��E�����瀚���i<�|܋3k�h��C͙>8Ѓ���PZh>�B:iu{�g�% ӈ�#�I�4�_}�����3���8��ҵ��ǫ(��E>a7Kd��N��i>��cX�r���}X�(Os�\��{���lH�zA�	;Z��L�šE_＝�Ma�;����n�ʦvx��o�űD�
w�i�Ǟ`ԁ�vw����}�JЁ�P�ջ�S�$����:��S��̪�����[ ����5���{qkq)�Pܡ�kJpww)Z�%-��ݝ�,����{�o�f�@&���=g�yvՇ��ً�ӡ�A>:.��\i-ч�������6�~�>�|#��B�u�{���e��u��~a[�������X�Kpmwi�P@�<�_=5]����T���%�Z%�h'a��+Sk{,�t�>��z21�q��5]D���B�/&v����g�D�|U7\R,�S������|���';��
�R"�{8 �z��4���z�~j��B�^�-ϊ�f����r�g+� :�NL鱸�G��h�q)ܳ���k,��m�C󂧺������mҏ�P�`Ņ�m @-�q�T;@k��P��B����u�O� ��/�#���%@ɻ:ߖ]+Y�b @��£�
Tc��Ƹ%́�q�r7�h?����e�:�dP�7ֵ�u���{��Ġ����:��OҤO�$}d���-GF��]�u���R@�W�����wZ��PB�3F�m�?$&��^�"=��* ��?��!�ġ� /�,T����:���&���:Ǜ���]� {Lç���@_�a���P[&�쨳IQ!iȸ��?=!��ݪ�eJ�n4����?J 'YY����_<Yxb�bvSu3��MW!�:�]�W��X�[VP�E=\��f\.(n�o�+iMdy��F����X(�a+ÑU_x˔oR�f2�EAj�%�<UH�Ǔ_!o��$;�����Zi~0����'� p��%0�X�'-2jo�_�&M~4�#ʢK�o���L҇#y׻�Kx1u-Ͻ��I��1�^n��mt���6�solQ^!���WS_+n$���T���|%6�)'�f�:b.!�q�2�ٰ/;>;��Z3S�~��3a���M�b�����xLV���#%���ZD\O6mmm�+;=�N͞�*�L�e��K�oc�a�Q&�]���n�����N�L#|����p��beh���)�7I봅��g�;^��QB�K�a=N��}�}c��n����!5[�>YMw$�@T)�~M��Ǔ��t{W%��&5<o\V�;?Op��˱lFC_^V����bk���)�o�Yi��������a�ҭ[���6�y]��VL@d~��4'�h��\���4 ˮ������f��k��*� (rI���ș�H[?4�%�k�.b�q��9@�,�$$Db�Ͷ����S���c���?���x�F�B�4hs��[��b��c��fA<lZe�]D�s� N%*����\��a���3��-2�O&x����F�bj��XbA�{�ի������G�c�}�O��(�J�F*��=�������^�q��毋����:j4�m�߼�/=����w�/1�w�
��7�J�`[��b�8݊���\v<pW1G�\�E��o�`�v�eA_����L[�h�8{�W�p��?�pt���d���@�3�'@a
�5���<��	1d6.F�&ԨMYt|��ס�5y��6��<�Kͣ������+mF��&$֖s�~�?Tl�u�͘ޅ�U��dj�ߨQ��v�T�{վ��;�`J[�;!3"nB@� ����E��f��U��G�AA!�j/�Ȍ�f�5-�g�n�"}Cң��7-�R�/?(��/UfgcUt��,V��}���?h��~y�����&�
�qC�2�4�9�~t&5.߹1�q�%ϨLY]�����$��p!�wc��Ǉ��+���U#pA���Ô{�2g�0(?U=����ވ��4x�[�t��<�s����v�,حLH�s<��vv���;�GM1�晭��	���#�0H_�Lj�ޖ}T��`S[�	�\���~�6���_8������R��	Q��f�Z��Q�/d��1����7�}�-�\/K���$
x�T�=���i��ϧ;�Y�y�e��򰆽f�W
M�q��;�_V?�'���q|S�F=9����X򾇺ެ�Pzi]����:)��~�_3�#�q�fX�5����� �U�k�����*�N͂�d�H�#����H���K��&�I�����+��W9N�W�
��ڻ$m��6
T�����t_�K�V;m˔��3OV�?�#�y��-	җ�c�-q>���8%[�5����հ5�񦕷���Ŧ�@���[�?0�呴T	���)�d[�E����NE��Yz9�_k(���m�^�*�@$�҃����s*K�ʁ��³M+K�Ll�R8�3�W�~��}�X�G��k|C��mAq��5���@)4�[L��U&�z��#F��aJ=ת�L��병O	:�[�8]�m��Ǹ��f;����ϪY�nN����ݵ������-)�H���������-;,2�\�w1�YJGG'7B�,g�[�_�{�D��YT�#���<飂��H�Wu�N������z�`kRO^(�`g�#��6� ��\o�]�ջ-
�k(Ǹ��=�-1H���\G~��*����+C�{�W3m
��#�\N��C��t�[�U�1<)$3�f����\��y%Ve�絫�N�H���OW�J�6��izf�x��V;o�/� ����|nl�7_+^׬��n����)�ՃW��8򥏂�ҍiE0��`#	�غ�^k��a7���	{��=n"�����nK/m0����k�^�!q��[7�)J�& /F����TF�ղ��p#n1_�Ga���h�2̃]�b�\)ac�m�Śh�Z����H�@���G�beת:��Շ�@U�)X�x�YUF*����Eh��B밶=���=�(�N�E�������L-!Td
c�5V͞Yg�3��@�|Ar����o�7����uy�����R(��^$1��K����~����˥�:R��EUv�ǉ!3Z�����9}��7�>�Z�FR��s��s�C)#���~�m闆{]Eq;�A1���z�;n�Q���b2���A�PV+���/�͏N.�Ə�o4�OJ0Q{�W�	��/6��]�5�C�t����,V�2�x88�1B��0}��Y���z���P;������Kp�w�D�_v0g<���})��Gv`�YvXT�HL����u�#��$'"؊K���C������=� s��?�;U��Vّ�|���m�����{y�~<�k�S��b�*��f��-`
Y!\�gq!������F���BTID��Q\3j�;���Ⲫ>���߆0�7X풞[=�7ܴ��!�zRsF����_өw�V|��Y����Zʂ��D��Vg�N�yHM�g�ʡ�#޺czԪ���*tg��'�_)�pQ\C=��K� ;�zъB��j`D��R�^D:E7r�R-q��K�}a��ՋA��q��vV`�<3��ǩ ۷��I��G�����b�����q�17�]��a�p���qlVW��/ED�x�ڴC�p�sn���2���`85��g�p�6ᴏ4; ��[��C.�w�v�
��Y�QtQD�T6���@�2��Cy�@�e��$JGn���)~�ἕ�=���p㸭�Iq����M1��E��CGۄ����M�g���蝡\ ��5"�}i<�R�9��[�nHĂH}���1���{���FiYe��a�M�Nf�CꎓC#&b��z�&ܡ��šZ�'|I��6����L\�Yd>L@|v���x+��xN��Ɩ��}�kOW�h��d�> �׿�ϸ<�4��8�=�'�n�|���	$`/��z*v��m���#��O.��a�E$$R�v(X�#i~tz��Z_�8pF�I�e��D�N�#G��{9�Nת�\s�&߄S�<��r�R�����}�`Z<�nò�2]���#��|>԰;Z�哮�T�R!~ʭ�'��x�Yԧ?2Ɋ��8^o`(�,hz����ƾ��w�NsF���,�7q៖cS�Y{���� :qoٟ�4<���8�D>Б�U�Q�����H��:g^R������"����)�3�r�wԙ�k�/��0�����0̮���g#팱�-�I�#�A��E-�C��xp�F|z�r�IBv�t� n'-���pc��&knYӊ-���)�4)�
7KM ��,nE�]�|���@(2�&��hH��p��x�O,��;�v3�}���|�e�G����Yr��?��n�}�br���C&b����\�����\H�	Uz���ӿa{5X�T�1�玮<��N!��\�ђ���P�;d`��G�J�Kj{�c6N=��C��`�,g�����B����[�B�f]�ն1�̑�z���˶&2��Q��!K�������⛿$�\�0������8��Ń����P{���I<��|R�"��R�� �^�>��
��qgnT��a������[Q���l>�6�� }��u{�.Ζ��m76����kvJ�;(�QWzg8� �""�F=���云���^ZQ~"K�/��	���d@���
�QGX_^e�`#1�BL5��_�ho��M��d6k�z�J�	&��N�o��eƭ���$���i�'�t캊,�D[�� �V�:*�T)J��%�uR����sP��j��-d\���t涞 �2;ӏ�������9�����u�Vv�^� ��}��R��Ŷ�����"�|��g�;V�9�ȧ?�+�N�r(agL�ǘ�A�+cO�\�R�h�����6Em�������c�K ��Γ�7�LKY(E��z�9�%�]~��G��j�w۫X���k嵺xc\\U���ى�����z��P�c��)b2�N�Z�zN�-u2��A�m�|���Mn�݈[��1����r� ������$���MFOꒄI���U��+NS�,0��N�ER�s<��4�5���G�)__�E�	C�>4(��e�!(�_�O�7�DG��$��>���|$4.�q�=�^�w�Wl��j�$���	�9�?xUk)�8�t���0Z��BwN����'�P�GOuc#vvۅB�M2���I���D�1����%qv�-$�&��ӝ�9�?�I�N{n�U��3T���ǈ?�&>^�d�En&�Ϗ�c�Fd	#k���덴Y�w.��A_m5C?�%@8U(ϐ�c%%:���ٰr<���9{�ЪSF���)6���<C�PΫ59�3��w�b�f",8�	�k�ǉ_�
#k�CaӤ�c�&�GP�{C%����������ڔ���쉚�ĦgR
�̽���h����P�7��a�,X��/f��'w(,�Q�_�
B�	����v���MY�j䘙�_�``��N$�Ig�2m�ǖ�@�B�)��|z%K}��70�?���H����9P^��zI��І#����{�#v���vE+���R�8z��sxff,\�dco��z9򧐷k7�&������Z�N�JWK���?�y����4���8�HC琚FԫD|3el����d`Ѫ��1���tw������R�����l��*�s��]L��� �'c�� ��y|M�%��B�Zߢ,w��%'�à\��߶%}�O*7H�J^_~� �@�x�^eɗB�	j ���A������{�{yn��L,N�X����F�{M�%$�k%\��kx��9��<[�>��5�8OW�,��k�cyܥ�տ�*i�����w�۷Ǟ���pO��G��DR6ז�~�����Jl����5t�"h�����=g�1�Ỳ��$�.�����WYMm��]�n{��_�ǅR��?��,Q_GbL��JO����]�+n���V]�L��r_����b�ŕ<f� ,!�dǏ<t'uV���ڡo1�ߕ8��ё���L����Żk'^�*����m�߾*D�c�3�
x1y8L�M��MH �E�=�l)Q�ż�Q��R�b�vL��(Y�d����7�T#֒:�h����9�8�[.*98ir,am
��4U)r�)1`�"HL�u���[k�K���%���w����o������Ff���,���ʻ��{�Pu*�d/��g_�n��@ه[�;��,�gC��K��"��Y�U�vu9F�ʵ�~t�4/��K�B!z�_i5/T�(�������U�G���(<[hÙ|�fw����Fh<ϿGv�]u�����Q3F���cЊ�������P~j4w�:�;`k1� �	��'�WY������(��C��n��f��t+�3����J�0��(,��C�rSe���s��.NV�/�/tU�>�P����禱�~ݱ�"�� Z��s�;�۰�f�|s�]����"�i=�J��5��@+�h���%�Z���ۦ:��}hPА��w��K%rj��,��2�(vjLzό�޶Z�lv_1�}�g���Yf����yߔ�6�Wt���!y��0*p�DV��w<��-�;�C�y��!�=;��4�䭞���&j�g�smޗ�r�zA���ףծ�BV��y��}�+r�l�9�ס����&2	2��*�;J7|ОJ�^�题�)�Ņ�����f�75�D�S��J��#��i\��8<o��0vO�b��D��a95d*Mj���Q8���/	ur2pm���o���;����bZq�K�Oʕ2�v
�;�}z��;y��@D#����z('����s�|��`��IR��z�k�m*��lTb����c^�?���K5�G����Q#��M���k�,�Ctt�0����K_�vTX��y-~�n uT��(Oȓ%Cn���{`�w�|HU�O�>�>�������l�uޑ���R�!ڤ�
�p[�*̋a�y��0���I**q	����ݪ�B��>]��J�Y&�\?̯��8x��ޫ���jH�Jcǳ���S��w���\t�%��Xv���	ؤ�Zk���h�� ��n��B�y-�l��G�R��fUH.�+���J:,�=�2A3��Q�y�Dag��;�a#	f��B�kn9�[L�fܝHڮ��6�Rn\����=����^]N��ON�z�	(���R�֚�x��>���m�� j��р�_:�����|ܹw�zTw��`d��٥�[�[�}p��bo�r�Ţ
A�� �_����+�{%��K�%I�>��z�'��>��H��L��vİ��O܀Y�]�� �]���d�~���A��uEԹI5�8o
ư�d3���@���X7̡F��!�s��3��#��[�h��p@����O$�"�zK�Y$�N&�A�%�[@�Pl*����1j�*V��ݿ�ݘ�b;�����;O�[�]�h�J�k������7�AT�:4b�uX%���<�,:�r����_���u��Ц.���+�ѳ��lq�T/��=����ߌ�꬚y�rȲ^�+�@�kUm;1;�?��4�
�G=�/Ub���i�I\�7��� �mx�
�O>Li}�A7Y�֕���V�z��x��.��$1i@J��#�S#�!�Ϳ�J�=����̹iJ҉e$�SI��_Bޒ����Wc�M��-Y�������?� [N�.Eu��B���}����3�[vl�7�ߞ���q��/��foVJ��q�|Up/�'�& ��nO�����{���2RF������\g���C�uB�����M�3���>3�|/��O�A˃��������B�>!������l��YA/f6�{�3t�k}P�}��x�n�G�/Șo�~�%�@���叇#lw����]��|�'�]�ln����p6�����a�3���,���8-�t������!�"���@TQ����Ԩ���uL���9R\D
�(i�ǣ�ܟj���Co�5ҁ��!,��l��������:���m�$�����v�r�,��������V+�hu����5�a�WY��&=ۖ!\����3��`�f�jX�Ϳ��9��w��H�T0�'9��*u�JX�z�^�����<��eХ�٫�مg�A���&x�4K�A�Ӽ�I��N%ۿ/��ĆS� �i��l�9=��
��gT\$��,m�G>����Li�Ù���՜hL�O���V�E~l�1�}�� _�i�B!�/��M�Ԇ'
�4�3�x]��C�evڲgdY8/MኞNu���f;7��d�k,%Ql��	����ӐA��ܲ�ё��4
����p:jQ���\=߼�c�8�q�Z\��	�;v�f��؀=W*ms�"�Z~�s�Uםro��*���1aeC���X�� ��E���&��sl�o|.�D�ʌi�5���v0�7�ϻ,�����.^�XyG�i�g?Ix�]�5��R�\<�:��ԃ��Z!�
\"|a�6TB��>�u..����|�,bS��A%�Zc>~`�.�j!�p0En��_�j�����,�:�w�w}�M�S}�D"�8�g2�	f��0Mz�T�s����b ��䫅��'f�?��
ِ�O�S3�Gm7��W��ߩ�� �G�O���dn�2�́ATF�W��ZחwH6y@���L�FUp�$�?K�~W6p ����P\SM����v�՜x[:��L-��8�2PW[���D˼(3���S�:� �3�R�y�l�9����1�����l����Jw}�ne�mS��	b��0Ŝ��܀D�.��T��w��c�,R#ng�VI37=��Dzi�gtʦ�`��$(���D���Q����A��68��i��-���9*ĵ_�ݩ�	~.�D���<`��A<�Z�[ً����S�{g�&~�c�Me��w��Fv>� a��7�4@lIi\\ ���X�SV��Ͷ�zN٣���,�̄6@��=e<ZVW�YF:%�AT��9�i�(�g�z$Fa�*M�qP{�\�@�$�j#��ô�oN>��IO��sk~,T샴?P���Z��k`<S��Yo�G����b�S�Yئ6MZ+�0=7���J�GYĹ���]g�y�
X��Vվ�]�4��j����m�t3����01(��|�~��d> ş�0�dp�;�OU��17�ă_��`���(��~���kμ��Ac)E�y�x�.}G?s�:-SEQ�`�_������Vө��Z���te������̝=�͋���8�����]����W�u{�ƻV����G����%f����2l��}�#ΣVbv9�󵈋;.�l9���E������%9NگC,:T���7�d^�w���k�*ͺ�#�5�����>�oLd��c4�'�՟J��D��|�$��4����̌V���+�F�B�4��q{�o���g���5悃ˋǩA�	�Dq���aF����b-c�b��/ʿ�p��g<J�\őe�9�C,���Kf#�������׎��d�h���E���suIh�X��|�pUlqqr�@�Y�A5��ʡ���T��I��{b��lC�S��m���g���.�c
�J�\�85�f�����q�h�iz
����]���L�W��/ҽ�ĘUsjN3�	 �E�j��v��ǲ�ҩ�-z����|�11n1�g?22���T�?j0�&!���L�fF
��8:���F$Y��������t�����੠���C�ړ1J�?���7=���Ό�L���9�$�"J�}ת��QD���ʻ8X��+���n�TW�r���0����:Cݺ�������P6F�hr�DU}Ԏ��b��k�Y�Z�*۟�r/A����}�	��[���c-���
7p �%+�aE:Ψi�_�s�I�r-��
h|�=�B�r,WƏ]d:5�8�����w׾�y����7r�����:�\�-�0�)��$��K����j�����<�)�t��<����<��y�M��Z� ���$���?I:bĚ~����^����.[��'�sq��=#�o�r�V|UV�ڤl-k���G�V�_�f�D�q���j�+W�蠮z��l=!&��L��@�?Q?��C�9K�����s��L����Y����<�Ǩ�wF���\y�f�(M媂՚K�B��3@�(=K�Ҝ���S��w�R"���uY���Aa��8�8�����*�a�d@+q����%lR>�	��������� l@���3!�B.�]6�Ԯ��eI3R�p���ޒޭ���  �9�x\N�H��x=�)�Hn��o����lc��u45C,���&��~��cqXw�z�zQ7h%�
��w�@C�Xo����7�~�C)y���Zq�]0�k�	l���������zN���Z�''��4r�$�\V�C�6���'����t��N'?���Y�+���C�ٌy'@�(�`�]����n�����$+T�`/PG���c��u9ca�^[CCc�0^�σ��韽X#�>c$c�Ȑ.�r�{u��c���b���|�ujTqMmMnELe:�@��p����i(Ԑ�9-�t��>YG�IJ*y�� ����K��"�6�(���!�IJn$�o����|�e��o]��ܟU>Hh����#�o9����g����un�vs�	i���C�i]���d��]�r�,v��~`f������u����G��|���
?'��k�=��������)�bHTI�. _OC�6E����Z뫵���4���}�,P=b�e�=:b��y* ��8�n�Щ3���s����x����yl��4������7_I 	[�2�����:mv����o|rm�����w�
�������Lv�c����	J�o��w.�)�w�=�5���Kk� )B�}�g������3Dw����
_��D5�q�)X q��H�َ؎z�2a�Ҍ����?�'��Scm��
�i��`�V)���}�lfOc�&$�5��a?e�h��!L+��MĿ7J���׻��ݐ�G�L=��2b��_���8��(9e ��b���f��ׂC[��0�r������v�M�X?�t2$_�y�"� You����s�\4��\���榿��8�fe���"�(�W��<=������ml�io�zI�9E4�"�|�	{��M��Az��1}�1��5��mơl�jv>�}�K��#�q�N���])�6�����D�� ?�����������=���EG����]�VX�p���*#ti�C����ON�N�}�٪���t�؜�`m���:٤���1�N�LT��a݇�e��s�IO�>���aQ��pC�-�w݌��-VS[����~+x[R� P���lix�&ix֦ř�B%5�l������e��cG~����z	����w�+���R�?� &��@s;X�w�1���c�
:7k��t/Me��Y����{�t�RQ���4np#6��ȳj��QU��xޢʆ�[�oa�qE{���_�M�O�P.�u3i����'���}b{G����b��n���Q|91�^W���I�I�����ާ}Dë8�'Q�J���Rd%!!�$�t���+"�ݎ�&��f#c������LV�*C��9�X�O�9���3�!�w����l7�bGW��:�R���y`�)����Q�]��$?���5>
r�����M��TN/8��+�����N��-���l��a��X1p�e�^G2E�5���t��ިT翇�-dh�v�K]���A���{�iǚћ��ޜ�0��c���ۭ���^�~��9���W&sC�ӎ�X��j pl�k��� 4��AO/�i�&�y&@S���	��� �	8be-��w�'Lԃ���M�~���H߲W4r�l̍������:����{ai,݋-�m{#-D��V	=�2	�Bv���M�_����M[	sCA�T�D��a>��A��}}�yI>����γ�%���S҂�i��	�z	�X���ςM)N���G��>�g�=ۜ���^E�h�oj.8����>�2˒������E>.P�|Ssh']�}����1�u"8r�����ʬ4M�4痃lam�tV�;�[�9���6橡����<�9�0��{�lfe��;����<ԥ\�&a�/����8��Ⱦqg�'\1Ps��`��)Fl�0-��&��;�$АE;B��΅$B�TY���#L�hiM1v,w�v][�{ ���6�Ö�B6����BV�PʅK�ۼ��W�sBH�'|ָQ�u]?��e���P��o���MZM�c�Ӥ��W;��E�xg�WI����r������Ɋ��Q�Y���))N��M���	"YB4�hi=a���JJ����O*��~���t����z�)d;��X�s ap_�U�UwG9+8����2߰c4�opru��D5���E���"���	`��ky�"��<ݴ�&����+:����\��ؐ��g��)�X949�����ڼ�IF�mWw
����N?�4�M��v�b���t�N����_��֭��W(4�z-#@����}���Q�Pt[�%��zڃ�8%ϵ^f�h����&��|:	[v�G�F�}���XG&.lI�0�R\G�f�{�}2�_�߾}�Y�3b<$A�2�p��H8wXi�˄d�9���N�K�~,ϻ$�mw�Q���~h�ӣ���-���N
tƴ�_^��������?���^���U�y�r{2���=�a���r��qO8�|����� ���a����o�!����7�J���{ay�T���Š�||W����F����4r�2�)�{־����"姯��:+���!���~ E��-�-�7Yr�ʧ���F����%9�ϵ��Ɏl%�B�ٷVu�ƽ1]��T�$R�Ĉ��m;|�/o��>�4���T�	z�|��RXX(�#�i�ьF��t���B���"�k���`��۱��u!ҕƳ����FP,��?���ܫu���.���|��+eJӈ��&�A���v���,i>=�e������O���i�Em*�^�hMV!�%�4g>;�!�x�*s$�Fȓ��[ʁ�bq�K�������� �UQ~�a��\L�$����~лSM��)g�R�����y�H�BX
��3|%�!���x\P����(Y*Wr���#8�xУ�#GKvc,KvRH=�J����(���J7
/���v�'����M�p���Dyp�sI����V�gQT��H�¨���ԣ��y�[�/:�h����	o7ܾS
S׋��b-�t{fQJ�"��W]&%v=a�U�2�ý�e�,3)�C�i��A��]�0^6�M���*�]�E��������;ڽ6���]���r6v��{9���Xh@�>�5���Jb̕7 a���J?ͮ,�%ē{���Q%�x�!�x��?G��*����{�Y�^�ՖJ�XpBg��f���pa@�D��9��RB�KE�V/��D�!(tJ��nQ;��
s1 ����-�B��+��#�8�p��6�"F������aQ��7�#{i�R�G<�ixa��{T$Β��J��"��0쳔H���y�y-��E���!	f�?�9ԓ9�����3}���󯔍�G��P(����q,}�p�
I���9�n#�N�]TdO��_�z�v->z+�k̔�ofTl�da(�UƉ���Hwc6$T��g�R���t����T�����ow����ߦ�*,���\����{��!��r��p�^�,.
����R�bk��� @�WL���:��Ǹz�鐷�Q�:�����7&91~9l��v���Umm���M�~(�� I�V�-�#V��B��䥖<�'n� ����NA����m~�J�0B���p���`}zRUmq�M�s2~a��8rUT�r�/�c�T"���k�<�l�R�]���y=��23k�aYGo:ƾ�TT�s��Ė�Q�/H����iV3U�ᘘ�f���1nbbAo�A�� Gz������W[������#1�V�� �gٔu�e����I=����2fm��8
a5�4d�����6 mR)��_[�:4��<�qI:�o���Jlb��uk�k[��0�J��4%�����?@nM;u��x�%砩�M�p�.bu�q-GS�r��������D�g��i���f��^z5������3��O��\��yb���w_�;�Aٷ���ӓи��`T��A��}���G�$�&���u;ݿ:1Z��2�`�?$+��C�f�_�H��4�'�)��"2�b� 3��`:y��R���;p�Se��q~L��%qۆ���w�&L5�1'J��n�u?z��]RTV���7K��]z�Fg�IoyQM��'*���?����Rȏs��n��U:�>�x���*Y��ъr.��2��g/�Ύ"�Hl��e�Zp{��@!_��sP['kI���q"~�c�꽥;fLV���4Q	�S�.E�wq_՗��߀�R��qY���8z{p����kc�#��ԋ8�lF�d��Ǫ}�FW7�O��m����-$����7��U���I9(@=K�����܀�&�0n�����s��t޹'J�A`U���l$[��<^:��)2Ǐ���~�A,A遁��I��p⩈"��4[��F���g3M]>���H����sf��6.�%z0�`���y�'��"E�B|��� �����@���{�/�@59!u��_��)�C�y.y���zY�xO|e�����P��+��	E������Q��C���%ũGtU, 0w[^^^dd�?��Ӷ/�)�l/#L�".)iF��@�vۗ}Ƈ-M"U��p6��x�g�;���̻ھW���o�^�� ���e�T�8V���I<����vjy��,��~�e��ߤ�	��a	��6c�u~r�v��>��j���$Sm[��D�<�h:�hnwf�l����+u���k3q����a۝�r�E�8�� " ���+z#��y��}t��drP`���^ ��|���p�ij���a(����~
�s�f]$Zf»��R�a?Gbe�m������d9�mb�7:�`	1{�
���ge?�q��T�en�;6"����H��A�ڹ�E�a��O��6�6%-�Z�q���m�ʼ�����5h�8
�C!���6}�~~/�_�=^	�πږGo���cWBs��g�}x㚥bGw�p�{�kG�ϰ{����#%��&xiCG�QZR�o<�4p�z�߷�fPDs4}����\��p�}V���!�2��q&!������c�51a�{�^<��\P~)�;Z�\��T�;�7"��J$�����A'�uԚ���w��+������ ��T���Z�o��6k���V�m��a�.���Oe��*Gv(��m�;�NZ B{f�IL�M5
�K+���_CP��GYM/���Y���5�A�p��9�2���,C˕];H����sa��V;+��č5y�T�R2D<��9����Rֈ۳G{l�in�?��YYY`�J�(P�S<¾��������PFgE������p紉3���;gu%o�F��B� ѡ3�<�ٴ�f��iPم��]�#]���뱈.N��7L��uR�����?QH�͑g��faW0>��$M5N�����P��AQ�`��+��ΰ���s� ��]�}
������>�fFs+̮3��]�p&navz����|r��h��.��\����

�i��BLNګ�z�Zgf	ܰ��è�mѬ��6��&���rs{J�h�kT�9`��<3F��Y3��2����!��V`�;�T����2x��L��Q���f���ڴ�чn�!RN��w(K���`ܞ�%.�,�e���]�Ȥ֟i關q�_6��@��_���X�2���N��;�+f�S~Ȳ�E����g��؜<��sǐ�8�� �Q���i�Ii��	���)�U�4��(����-Va�7�yG���W����ĎS���<��Z�����j.��m<ߥX��O���d���.z0���չ��[���^~6��z	���Gm�s���V����6
.���Vd�@y�,\���g� 2�t�$�12��J��o�O_�7�4��\η�f!�6!�����c�6�u��^�Lgy�I3+(�	��P����-�Q��L
>�96�1K뼱AöEw2��L�\���t��A`��8�T0��PK�I������:�_bđ>�`�O�Wq�=Bhi�C����;i֨�"Lp�@Fn�q�P:��Z�����Uܬv���bw1�<��[�4��pFRLp�qd�G�y��ж�*��zH�ٺIn̚y3Q���i�֛�<ՏZ����p瀕�|j�B���1�z���8.��:n�Ȣ]߂yUX��ñ������l�u�[��61�j)����;�ST=����	;���w##sϬ,n.�/!���D3S�Ӎ�v��������$�4	�
��+bNG��D����+Z��a&�#�?2�.j�9��
5K���fA)�m��մ��b����O^�a�̈Ƨ�)����Ւ���أ\�͊�ݠ���L�}V/����R�����46�]i����%�;z ��(o��a�&\�И���hљPJ&�w^*<ĸ}�BRKKK!�����$���֗^7XY�rN���wY����Bحu�7 �!�w٠�t�K��.-Q���H3B�N�Qc�[��AD�0|�� ��F"�z-��£YL�5eE�É:�y8!|}iڻ����L�s�z�c�:Z���eAg擟v�޷u�����O_�v�}M)������w(P�X� ����
�X!�J��Z,�]��~���f��2�d��=��wם���`snڹ	�;�t�M���|G�pN�T<��U&QLY�Qn�2�9[�_v ���upበtC.���*��u����Ȗ̯X�B6��������V��\<v(�?|0�ܖ�r?emr�:����1��AR��8��ܩ���OVPo�Qg��~29��2�\!�l��	Pe�"�hn��у�ќ{q��稡;i�,�[�Y������+�� ���O����6z����Ӷ6�{�nٿ��K�gu�ӂ�?Q'~�N��3�"3�m'���o�t��(�b�!������ܑh�����^��5�6"���E-u�E�,c����+���P��3�f�����m��W+�$���M9�ݭ2.��T 5��>-V���|;=P/�l���(TG�Q3
�nl���E�6�Im�&H�!~��{�Dl���&~����(Gh�5���i�i��Lz�����%)W��q�k�C{��1mITkwjz���Ժ���̧�D�m�FmT���!g�6sMC!�DD��>�-��Ww8!�leVG�fLX�o��D%���+�C�o��p�LBJj|�ZX�AY����us���o�����צ�Ǯ`����_}E�����CGr촹.ς	���<��i
�kU1���x���1�����95y��@��7UF���N7g3 *w���C-crlX�گ�2��n������j�+Wz������qf����8����a���$$s�I;0��;ȶ�Cm	�+>��[�{���`o`�C�J��G�=?�+fd�[�T/Х��sݘ��ZʣV�f�5�*`&������ԴC6���p�A��2�hE�)l��@���3ؘ�ׄ�Y�~�_�_����U����M�Zsek���&w���:�/��N���x�bf>�Oʹ��^�+���?d�]p��=γ���)��-�ǫY��=�5��gf�Xҗ��Jzo���b�t�~=����I��]_%��!d�� �{�i.dF�%��E:w��;=I	�8�ngh���_��D��:#�k���@n�ū��;W�Z��΋)��3�Zm��[.�3^p��۾י|��~�ɣ�hQ��u��8�h��><��&�r:��{ؘ����JL��_�R�9�蟇��Os�"ȈOk#"Z�"�����	Z�H��]�N��#ve�Է���j1�-�.��6V����>(g�.��#�׀�$�Yi\j.��:	��Ϲ�[y�Q4�[���*9�{�(�Z�B3S&���H��b`B]U H��t�mL���B��Xt�T��'��UҒ7\0�5Gzb_	�dud���ך#��6i��	jQ��=�?��������R זOOG�������������l�����c�@���v�+��U���,�m:i�y���q)�#A���1��hɞ�w�Z�z���f��~u	D�m=���N'h��-ى��a����h�����=�P/Y�z�-+�T;Wv��)�g��,��]��
�#S���6h:B��zKwK�9��YGc��|�;��:&���9������!M��{́޽ő��c{${r�3ߧY$ۓ��sV[P�K��Sݖf�W=��Ô���6{V���m���O�*U��Z[r���e��%�Lzyd���r"W���.$8F��q�ٟ����K�wY�ҙ.O���x ��)��V[�/�>��wF�S�?ASV�*<�,�6���ӝ�^�9�;M�Kľvf����H������Iݹj�o��[�~�5l���u������u��mݛb���_���kFIU<�r1b�a�<`��4�����|��j�<U�VB�J8Ҽ�3�dH�U��h1�4F�zӥ���0��B I��!�h��@��6�H5Ԙ����->�*���,]����h_�u:�bu��f��}Tx�oJZ�&J'�{���ӱ��������2y���?�N���ԋV׭���#�Fj�@U���]�+a��\V���0��IɌ��$�ѳ>��@��
Nz�Nׄ��MY]�3%�ߴ�i·hA�fFFK�,�Dd���K7do1��?B�@�Ԏ��}Tx�<����`����f˟�dq!!���!7���\�X��q����3-��m��hA�Z~B�IaR�fR"ҋ2/��T?��)+�b�|����k�>��T;r���lv�B��/���`�����gk��
>��lg<e�Cr��D�V��5��E=��H;��Æ�ME,�%Ӯ�K�@�rmC,S��M��T��U���L���S�N'��㭗��&H?ܸbF�.עqz����nd�t����X�]˭.v���H ��
`1[��t-X��,p�R����K��mc�����h�(�����qZ�������_�0�@����t���rt>�LNL�f���Y����"�i�=��8怴��
�������A�Ԏ|�m�˦}���_� �X�Z���Pf����֦zi�qL=��6�<Bf�	#H��߸?(�����3VC#��~����W�S�4c�_���r��"l7c� w� �)���B��6]��B�O4bzi �4�^V��;90�~^nkb���2R�~%��b��r)��I	ڌ�os�J���M���G��d�/�T��RR�b$���
���e'�爼~��(��)&@��H��"�R�t3E.(��$�-^�&�f�����b׸��9��S�����OE�;�7��������dP��G^Wb��;>>lP]�U'	A�q����߰*�3,o7�C�ۗ��26�$�%��k�9I���?�a�2v�)}������}�������땀N���bG�}�
���`�A9���.D0)[� ���~)�X�/�&Y�s ?�~��+�X����$�)";*�#���lW��7�`�y�:i��U^I9,�S��<�ɒ�p�/^�Xb��'��ns|]jO�0&�$ ��eۖݻ��4���D:��� ����u�u���B�؏����\��^��%#Sdb��Zo#0�G"��k0>�Ƿ�,w��0���s��c����fסdpc�/"����\9�6_T	E���q��3�gU(k����"ϮV���YJZ���2sT�C�|��[�����x���xց�� A�!�y�����9��LFԚ$Kp6.�ޡ$����*y�)R�znIێ��;��ib��v�~�9^t���{�Os3��D�*�$��)#�T`���sF$.�#Z�zW�H����8	=ذ�)�_ �K�?�n���l���\s��r�.c)H��Rﲧa���^��2ig���'��f�ң����e'�;P�їd����v�_���Wv��+���6
�S��&�Q������?�4:P�ΑIEl�	����>X��վ������=��Y�4A/��63����3�*9��C���\�� D �#8f$����
��޵w��\�ztG�)�e ���f�M�P<]*���:���8���m��̊�o��O����1�K��O�q-��i��#U��S����p!���_�Ut�/����̍�"h��!������}p��}�b�Z��'���d)��@��n<3
�~̟�3�ʲ�j}��Uo:�[6�����l��6�O����vB���H!�w�5��s�΃@���.��!t��ￃ<;0��l՝*Wt�S7u|�1�:l.�́axd#�ɢ�&�c�{��?����7�6`V��㚑�����o��8V��q6�W?`��eWd���P���꛺Q�Oħ�����q�0�� T�k�8��{xMk`�@3H������C��ͷ�}���
��-"����CJX����R��X��n����?��mo�b��8��#k+ip~~����}��K�a�QE�s>!�<A��*�_�F�{S��N�9�x��ÿ��s�4��rp/ԙ	ˎ����Zj+�i�Z�����ڒbJb��\&ݜ���X:��agG�E=ݗ���z��f<��~�I���mc~�"��������ZIh��%�w�zp�_�>t��K�����A��۪��T7���ʹ@�������cF�nݥ��d�^%�I�K�l^�|��D��d�U�BZ��:�|�[w�A���Y"�q�H�5Kr�����t2���c���pQ�2_��n�턘7#ݶruu(��v�ǉ����o_P����%��D���:n�8�p_2(k*��w\�I��_E��A' �矛D�:y����+b9��[�gLFG�U�4S���!�n��M���A�SY�����KǚO?���ki`���s���Xg�@C�������8��Up)E�ӵrhp�J9A�4�����_t��6�M+{'{����o���&Ã����6;�X���5��I
�c����ik/�ȓXdY��I����8���Cz����� ~�Ҽ�Q�N6��j(�D�~ن�4��Ґ7_O�/��{��ap��\-v�=4ۚ4��Z%�}�`Jw�����\�W�s~��S�frٌ=��Zn��q��.���6���b���QRn�?�p��>�0n�����bj�q~�
S��^1���l=��D`s�����&x7�%ν.�
���4y|N~!��4�� ��M��QeoQ�p~�{Alk���	�MX 1��v��`���H>�G������yԅA��zgpu�b!��b��22Ys�.q,LH	��@��QG�0E�Pt^�ӵ�k�=DN�,��T���恑���T�z7�~�}F"EP!.�O2��TƕHW7k����1-�c���~W�A��N]�;w<A3�	$�)�
 H����#�1��������bR���~33�4C7)��}[��_.. ,�D�^@� n������'�<�u�������߮^�$7U�Ys���ϐ��3�[���=�i6=������l�F��)BPWZ���~)�����?l��%�4�|�V�I o�9ߢV���b�
��i��3J5�^���KZy����HV@����-n��3��q�p�±����7g�CW�ޔ5J�Dg?�o�7ۤ�_����.(�����Oګ��K�a@F�+b�tI��L�z�G'��i#4�xkύ�E�R�ã�N5y]VG��J�N��S�_ ���a���7a�*΋3C��,J�ښR,�s�y�]@0��o��_�G��Tp�:���3����׾�&���[�wr�T�: ���-��S��_c�1�ҷ�o�<h����+�9�Q�r�PP�B�9���S&�ﻚ�&cr�-��O@K遬��j9O�=[?�j��	���q���3�eTgk�Ii�kl7��hg�q)~�y4�����i7�HS$4&_�C}�����F�w�*Vș9�e��{Z��V�������^g�%��i�&�Ǣ\��s�E����������%'�gsJ�5�/��z������5&aIQ1���>�5UP_݈Wj���o������r�	��t~������Ҽ���c^��b.�GU)�$�͛Sa�r7(�K�n[���'s�o�_�w�F�L�`������h���V%�!���y��?�I"�\,���{T��Rz9�V��o�-��q��t=��&��jm��k���&�H�<۷Mt�lA�q`����y���p����\�z���3����\������l���w�Ŕ{�RtmBV�ƾ���k�ə���:P�2�A�~J:j}_��d�;��������>�'�A �h�bss�q	�~�2k���2���]��3W[�n��<��z/���0�d1a���|h�]ck�o���y��-�K��`������&�J0�
�5!T#�)��9y��N��ɭC�dHs𻥩'�GL�Jc�����ip��cB�\(��#q#�mi��J!�qԻ�hW������U�0C��o�N�����y�o��O4�},ú>�d�Ȃ���z�yQ��L�<9��oK]>j9o"�rm����EJ�O�ޝ11����oe�����`u�OaBY��us���văl^�1a,
�<h��k���y|yDA~���%�ON��n:�ݵ+��mܨ��|fȃ�K�s���f�֘N�MY��%]$!W�?,BÜ���z+�feMm=��)z���?W�%<X߭�����%���gCC��;�wT�ؾl.0��P��k+<�l�PY����P� ��Z�G�7I�<�[�:�`�t���5c�}�4c?U������2���sD���㕪�[�QC}ݨ�3�G^R{��ͫ���r�֗�X?2���[�#8��M�뉞ku�k�wܑT�Ft�]��vmJ>~�J
v��^�<Y�IԄև�̪�H���ɟ��ƫt<6�����5ײe����3A0PW�F�Ҝ��2�^Dq)Tt����eI�X�(#g@<�m���QR11m[�N>�7�BJ��n�"E��T<m��c���S�Qb9`����O��LM�I��I�A���0�Q�����i�/��k{��2j������6X�Et)�kW|a�Ý�������{�ڔ2B����#���N�8Bv�n (�i�_�����Q2ޟgq��HB����պ��'dD��U���'c䃙�a�=��򺅘sª�2ƌ�M��h��Q�s�Q���-��:#���sE�����q��O%.�Y֧~l��1�0�#=���WD�{�v�::�m�>:*�sIm�&%�!��-�%��YN�!�t�����H�mWTeqr4[�K�Rq���WL�=x�VV�6	t4����n
��[l��Fv8z�Q�?���5�M_�=���%�Wr��҆k����#�l�(�Y	.�ӷ��1`!���b�H/��e�m��/%��֧>���L��E?�W�,ζ��7�BS]�4L8�Xtٚ�,,�T6�q>`�w�n�HB�����ș�/]��[��w=�-�~N��ri�#o��q�]�e���E>��(�<���^��c|��k��w!ۿ��;T��s:i���5i�l�/���ɺ��u,�xu-����<M�2�z�ɏ�%��Y��7�P%�>�ӑ��B[U��9�����`V�3s�$s�o���w#�$䣐�,�׻6��Y'\!� ϊO�-���y>��w�U���G�D��[]�_RK
�)�ӥf�f�FP�,�?���6��x,�܈ <��&4�E�k7��jx�.k�@�&��#����ՙ<&M-��w�cK�>�3Y����`w�6C>}�a����ugv�.`����P��w}�)�˃O�Bv�tͬ��������_�ɺ'����A�:��o�y��NeE���T݀�S5X��ƻ����iƾfu~�@�����<u������2IKK��_���{mB{�6��x���~��k�
�� ��5�.<r;=��&��:Y��9��I�x����CnR+E�m�61���������%��\�v�������U1s� P���8U�[��q������~/�������Njdo�g��8<��SB�r���{��@[���� ����?���j�X�i��z�kt�_������
���teC�#[�7S���1��O�|�S&x1jm�c�yZ������Q��B�3 G�OA;�����X�$�hJ����T� �z�V&��9���Q8&��1�:P�p���Z�<v��t>�7��]ko�'�RjBi�u<�E����l���
٦B�Ts
���^=�=jM��v�����;zbd+�lJ]����s~�I��~.V�k��+�Ԛ�l7�\3����.c�<�9���0x���qŜ�����x:/�r+���%y�.���ￕ&�R�ؒrr��,,�QѨںڒZ|���U���c<�ؚ���З8�^�e�[��p�Ѷ���5fE�e�����卜N!3�t!vQ�`pW �֏����S�,��Ʌ%������h�KK�_h�R1�ejVo�<O���t߹\/yX�M���loE[�s����R:�n2�5����
�Ey*�.3=��y��Yjj��diT�[��"pQ��3���6�z��T^�RG�E&��d��N�V���j�è�Jo���bs� 1�7~��7�ـ�69N2��n}�ʠP�H$/�ī���ɽ�h9<P��n|���ooK�V���	Yuݹ�V�o��LE� e0n�7�18�k�*Gp�t��PA>?\y���m�9�Fl㑗�C)���q��"2t��Xb���i�=|ﶶə�P��#I�I*81������N�����}��F29�t�W �bb6�vr�>o��> /�j����!݇���]�].�HBw?{�.�^����0�?�9������Zym\�ڳ�0A��+�hȠk�����j���M<�[l�i� �G�<ې� ��_	���xT5��H�X������0؅)��}I%�yGKK��T���/�R��,)f��1�e�r|f���L�IC.~I�$k��O�����rG�����$D-���B�h(�Dml������R�=X�eqab=���[z���n���}��pX�+~��x��������j'/D�q��R��7f��M��)���G��f�g�s�ޅ���=۷}��G�	}_~��`��BZ����t��,?v�ɷ1`BR�.Nsg�˘r� )����~����3}��_տ�vj�E��Vw�и�^�z��FI��:�0zO�,�z"u���hn$�ĿQ ��cQ�+a[[������}�[J����H������р�c���{�ِy�3�����L����`٢���I��)�ZѶ-z��o����^����ң��·
��Dc�e�TD��j�Q-��H-�؏��j����Qo@u���'W��D�k��Pj�R԰�������a����(�C��Ad��w���j��xQH�U��RDj��*@�\J�tn�}2fD���WXI���+�>^K8��9Ҙ�5̫bb�@dK�%���A��I{��!�h��8��ډd|�dۉ�%����$H�nԵ6Y���m:k�:r������ى`��s~�Dy�W*2�Y��U?"C�B����+m!Q��nnn���b�w�e��Eߛ��[���ܽ���	D|9=$6���~�������+OG{3a6�9 �ؿ�s���<�:���1yvs۠�䁈a1�4�����a0Tb+�D��	·� ģ���}U�#����éA���r؄�O´Ԥ\]y^:�v��r�py_k3IK&��E���:V"߁f:�%���z�LD�Uj&M���6�>���f�k��nsU�Ƭ��Y�� y�@�#������%֣*��6�vB�����N�֚�+��������9��� �F�-P�� �@O�0��ӓ��Cqa��H�A�ȄM�]�E�RO��[>��k�R���f�Z5<��p��B4T��IH<`Pe��{G �vDX�jwEA~��{�ܑ�J_u�;���0X2�>��X��D(^A^(�ݩ��闫FF���Y�M��x��?�~��	łY�kD"���y钥Jl��\���)B
LG2��)��'0^��j�x�G8P��Ҧ}28v����1�{A����IFJ�T���@BBZ۹�^���4���� ���p"ŵ� -��T����!����~�>|47UI,�m	�C����|���$� G�m���>��;��XF��S*�������&�У��� ������]���!�?����EoVC<w�<Z��5���ns/��г�����*+��{TM���K�+�z&�����'h�l���:����&���_u�1;���2����Q�}2�@C5@瞴���k쨨���),�C��:�~qqaz2��;��� ԙ546Z�}%��m����mhj2�.Q�m��5���@��c�0R�+$�W�� 2ۏ��oн ���`�\��|9�BOW�t�m�ԭ�EG|�jʔ
�X�M+�� ����f���^�ڬ�e��W���L�+��XR��zH�h�=�'5c�{9�����A��[���E{
9�"8�a�/���.�̨�*�؏f���H��,,���=:)�:��KR�̩+��]7�SVs�5ɬ�����W���;�Oe�#M���W�-��k���BLPo9��{Y'Xq��8K�;�-��pZ[O��8�^�����-�|����	ψ���H�~�ֿ�ϙ_���!�r�{�6 eˁ�0`�I�к!������թl�h��������3�5���+�����s�������Q7Sm/U}y��t�Q��UPh��[b}�u�����w[e✝wTj�"��Gߢ--K�9^K�V{O{�C�>/C%���v&A��.�R�$ta�a.��Xr���
j�Z"����(�j�������k���i��֥*Z[[[/G��X��CD	�~u(��s},��*a͚��G$L�7��Ԃ[�l>;g(`��bw����֔����y,r`����1���\����y���<�ix��M����+��nŮ��d����Y��+����ى!�h>�Ǽ.���@�]��g|NN�K��"�UTa�6�AhE��
#�hDe #K��}G�t5d�}���R��[�Q݁����G�1c(a$l�9�ts1/�����l�[��||w^�'����p���p((�]��,x, �99�hk"}�U'@����t��&(�E���ϖ��88��uk2.Կ��:,baa��:���� R]����"�����Q���n:� �t"ZՉt�'C2ЇP��ֶ�8�G!��R��lmp[O��� ������o݃i�A��:{�6��cҤ������P���nӐ|۽��Rot; �*�@I��Ҥ��!ߓ�j4�o5vKQYd�M��,W��ӓD]E�7���}�-�����#b.��g�4�).�M��:�FB�D���±�Q������6��ѳ`q�QPJ'�~~J�{�=��3�b"�=nLs���<8.i)�DO�9� ݎ
er�]>��[�,�B��#��o�[.w��;�����$�ߟ�f��E5�a�G�-�m���)��~����}?�|IWz$j={�_VZ��Z9����N��5o>���@��]&��6q�%$�;��vt�uIc���d��0��cg�x�#�|����mh���z�bd�Uo�F&����,�LČ�P�`k5���SmG���ҟ՝Phjz:��d�/���0����t$�����KY{049��_aޒ�'�'�xOw4��Ki������`����r iU�&�+G1W����U����� �+�e�܋���cQ	��Hb���.wG8�?�­5D.[�b�B���s��Ė�Ի����W�W��@퀖zk��N٠�o_(��g�(��g�{�3��A�6,��8V�8DA�\
��G���]<�]����	�p�\A�f��~������^����;��@��Zw@,Byhd����nt]	�IrugN��tS`C�x��gY��2,cbz�u�����ܳ�yKI�:x8�vg��V���'79�B(6�XI^upu�Ĩ Гk���>X`Bp��C�2�Á���K��5�����D]2�RM��u�J��<�1�f�aw�� �S���kg�'`_�nu&��e)�/�U���GH�iao�!-�&��_��)���h�q#��BgCl�	��
��@r<zy���Ef{L����ME�Ҹq�K�,�䞣w��]F^E�(�U�b�𤋮���Í`��`�����|��������&Я��0c��2��3����}*n���K���[��x��WРұ_4O@#��ӊz��S^�5 P�j��CD3=�;Cz���*�xߪVM4P���np�Bq��O�u��)/�)OT�f|�@�R���-Jv=�v#d�pW�� � %?/�VA�u�.����&�$�`��#D3�P��t��㊄��B�1�����́�K����y����/AaYș8;�<��[C���{|�uύ���x����l��r./��H.2�$M^���}�Ŝj��ٶ}�IYv�E:k7ϳ?⒱�)�id�~�������/���lm��`
z������q�} ��8���u�Y�o,}"4AU��*��Yn��,6��^ɩY"�^D�3�Q7W߄.���9.J��Fs6~��:j����UV���V���[+��ot��m:�W��M��<�E띉�b/�I�S;#�J�� ��\�B�<'�A�ir��Na�����煉l�K���ިפ`Ѓ�U%BvE���`,�8n�W��#
߻�RO��)��H���y���ђ]Z�t����n-��w��)2��W?��A��'����^�Df�����vh���P��K��λf`wЉ0ܵ�
�=Rts��2a�r�g6�ϓ5AB���6��N�	b��B����r�n����/7NMvH�@&}�lL_���(�
�v�-��2���L���]5̿bDV�]�_Q��с^Ŗ%X�	91J,I����Ә��_Ϳ,�X��*�![P鉒�t<���gy���|��Y�s���(a2jh���9( ������M]4A��B��s GuǗe$�~��ٟ����#�.��c�$Q�O��"��:e��ۍ��;�M'���+�+�wگ�yZ���&�|��X8�_䉼~��ް�v��xTn�3�[9hq6�̇��r���� '��X��I�L���W�!�SDJ?ck�	mS��\�r�[�z���(���eu����AFLr���k���[X=�q�0ø�c��H^�v3=^��<hĘ"*A����Y��_4��%y�)���L�*�q�m��}�n�+\�F�����Յ�|Y�k�(��n"�Q�Au'E�)�$ "w[W%�8u�����Xf������LIG�WM�/�#'Q�ۊ��)D�� ��\|�7�T�߬����r���L��>�,y�m�Bs���Z�L>k~l���oL݆�6�@�9�~���Bd�gu�q�l�c:���3�j�m�c�ms�QLKo�����'��&鹫��O��"�u��W7�ޒ
�3!��U����`P����$(�ԉx�򡨵
�mvN��:��͸;��~�~��@��W`���t��W
��.���E� �
&��G�������:���vG��u�U��P!Q�ޤ1M)!(��@���Ӱi�>Z����D|�_�Uݵ1�2���і5�&����]�}�+>�.ح9���:��N+�Ԍ����x����p���ʐE�7������P|�8;�\�=���0����	���Y�������3P��VÞN�k�N��K���F�W!zЈ��:8`U>^����|��9913�e���~t��%���R��J�|�] �u�P��ر{�������� �����C�in}mG��������y���/R�2�_��>},+���Q_�#������N���j���h�[LbI;����݃2�u�4Jo�nsʜϭ���ytk��q��g����7p�xU�,k�%'����R�%(^nJKy�	4�1}Y|HZ)WM����n����@.]Q�"2��Դ����=:�LI
�����^!z�~R�̟"V|���U�.grwv��8,X����?����ִN���[���$ʒ�H�yR׽�`53�����5�p�ӓ|7�s��z�m�����i��p�`�g�U�|Q��0�8�@�c'�F�o5����pWӑ?'��]hO�Tg�����1Ϯ?���0��޴~7�h|q[s����m'�p9�l|������k6fV�3����h�A�T�&)���`�	��f�ۣ��$�IcL����:0ȷ[e�Ź����0A� l٘;W���n� F���]Ȋ+�����<��v��Xw�R�J��SB��	R�s@K�]��'�~�T�H���]�Ϣv�d-C�.��j����j��k���}�_��Ү`G� dac!:��XTB�?�ţ�Uh3��9N�5D��=&��/������-}<�5�Zc<��9�*)a�v�_gQ�쁩�ǁ�#���icJ����$�"o~�����~=��̡����!<`cv`�z��?��"�X_U61^:��w/5�:��y��֊���tл�z��朊#oo�ɖ��86�\��0���V��C�wF޵С�D������yk52���:�����*��1	bB�S"h����zI�P[iO�����E�D���/(a���w��Ƭ�g��tl�Ӎ����Y���ϑzH:W��6T\}	"�Y_PR�����)�g{����AtA���U[W׼?ՖHScW������xU�.�	�<o���
I�ֈ��**��t�~-��8ώ�
���� ��Wf�c��n�4=��"���*XF�u����[�$����~��\j��!j���TLd���(��R2���΂�~��ɉX	�t1[_'�^(�P�M�Dރn�)܁�{�Cz���`�$Cm-��TW\�8�z�16��!�Ђ��Qv앸��"�W��,nn˝�A	��OClՌ6���XȺ�=4�q��x�i��ZΈ���:-���(H|}�*K��l�a؄��1�((�-e�~�7���%�	�:����@�Tc���8h�7���E�lXz�
���r�Y�8f��+1��n�O�$2D��~� �|�/��p��K�CJ21_�1����rs��^q
��Pj;����j`�_��닉�E�G�i%
hd�uƐ�	��H��蹜����-���Ⱦ���Ͻ�jW/�}��oNܙ3�N�7�ĥ�$o�,o>\>E2���[�Aq�0$3��Ǒ��1WZt�I̋�3K��|�>6]>��=���Cw��&^���ZT��?�H��Y"����S����]�7Jns�+��C�-�6A�'��FF��%�f�ݏÐ��P����W;T%���B4�:���Eo�'�_�?�.还��~����r�1(���ɻ?='�����dm�;���U�lY[�����m�?	1��G6~��*z��o�[�}���pq376��1Ŗ�ª����"��!M
X�E~D���Z�e)�y//j��/ו�i�U��ݲ�jH�Ռn����P8��M��ʪ����'�כ1��*1���A��=�4ڦ2���j�F�}02�7_g���u�����ii>(�rO���0�)ҽ����9�&k�fub�ڠ�8H���ᜅ�,���Аt���5����A�JNx4�J����)��r���Y1]���va���Fp��A�<	))ࠪy�A�6JG����w� ����rl�MlUVxx|�)]_p�?�U���!}���W�]~R���@�7a>�T;_zQ�Y�2��.�?�_��������Ø��z�&q/p��M�Z�h���tTP&0`�q�n�9�.|���� �:P�$�N9n:>���`v��0�W��B��Q�[Z�y�
k��y!Wf}u���8�馉s�
� } 1��ݽ=)y�c���"����EL�Z|�,XP.7~�Gy�q�gu9s���u���7#����H�-^�O�������s8�o��$��!f5��qyh,��a���W0�+��M��R���I���K���T��ddrKKb6���CE"i-�]B�0�4�B�/4�{,�E�P(��O�X�Y���Gya�	�U�nK�c��ۇ���,���I��ek��Զ���+�E�'�$$�G�����|��8���7�W���9�,�hi�䷥qh�HnӪWgs�>6,�ik��[d�,�cHNC�rG��z4�DTa���OX�S_(
j+��"=<]UD3K6��{�ַ�?ؘ���Uڃ<$b�2|�-"�6;��,�KW}#��C$�Ϋ[�0F���q��P���-'�{�)�NA�yE&ވ�V�b
��)���6��R�6t�<Utii�����Z�t�!�O��{��ق�����&c"����Z.t_8������aV7�GS�(��,fTo@<�l�Qz���K�����:�f�S�ӛ��jE����հ��1�㎈
�|� {�m2��,Q��4�H�0���xi��+�f��1cϣ,�GU�uڼ��� -�F�;<�I���7���v��Q�/�Tک堫٦î��#�q� CA,1�~�B����%�a�>����؍ ����'yT�[A��"p=���ewW�r+�I�6TR�
)Z'+���b�����K��q�8�
K,8�t�V�A>�wz:J��	�82�r��q��m_#hҙOA�����;��k�d��F�[8���
��޶����>)x� 3�]��ǿ���>�>�S	v������LN�П9�aV�	����:�̃`�%FW����4AGG����aO6��r�	$aџ��}۷h��NR:˵Qk+T������ފ�u����c�T�Z��Qt�0ij�l�w2vv�e�WėY¹�)��H������i� �3s����Hc��f9>�#
���A��/�L2�C���q,L�);�c̉����@GC;�E�����j,�����M7eU������6��}�m>�z�r ٛ��[�E1�a&<�?��:*�����S:��S�.I��隡�SD�AA��ia�!��!���{���5���ଳ�����s,���·�ArA�7A�?ҏ��k��F�X��T����'d�Þ��n����]]</SLL��Ŭ�$��o�&����i���[Wv�"�Q�d=K�
 ���/݂�1�ۼ:|[ǥ��W�v2u����u9Y��u���w=�vࡪ�W?^EU���'Yk-��\]��sw�Z�x�|�@�����;{Z':R��~?$?�JKKN����P�@u�޼+���k7b���#�h���OMV��g���}�viݧQ���@1Gl�0���-��ڮ���L�&;	_��p�nl?Y��-�]��/Fŗ�������s��OKio�U�;��Z}8�k�gn�ך~���DZ�h���j��*EHb

�u4I�c�&��׳�lmK]��gA|�+��BGG�ւ=r�9�GE������3;4E�f�ŕ��ۿ����1�ϑ��$����������_
!��&���Fh�Pq�R)�l0���Z�u�⽞pu��x 	UaN�ñ�WN�$rZN�:V��y �p�!�ig!�0���G��*���Δ�јe�ϞKp�͇/I�d�c;��	bEU��R{�C�kB5�Zx�Z:��ӌ��v�������-��.�V�B����"�u��9>a�zZl��{:�-��F��Ġ==���.������]�YI�?�����Djk�>'�@/��ʂ	v��/�����X��U
���;��I�0Zt6�}��w-�dq0���m���/�ϛ}ha�4sE�Eg���V_.$�4٦��_��*1[�=�o�Q��>���c��P.W����yj�2�NVv���b���Y�W�/"E<���L��&4p�w���|�L�Th=��!��C<�@ ?��4I)�i�r@�Ԋm�}��{��� ��f1 �d�$D�~����H�?&���,�$����Í�d4ùJ� #��-��E�?JNK�Wd�s�G!��ݫY�[ſ�Ԛ�����fP�LS�D|�}M/r*�Z�uw���v��X�ť�njW�Ly�Z̨����¸���紲4�ӑ�"�vg��|��e���L���Svb�߆W���WP��oT+��0rj�*kj��!����[�����A0�i��N�Z����;�^[��Gi�N��&雗�~�T�ߧ$�>\cz~l�lזy5_��w���	w��9��.S�x�$4�~E�Qa
�r>��h�4��܅�K�*^b��d�?8��Tֶ����d>���8�&��3�>��2W��vvj�Xp�!>ٌ-�oO���'���a%���10��AW��$ؓ[ �,����%��J7[t���c�YAi��f
+(�*��xr���6&C'�)nw�}^�������k�$��_2$�=�%U�������1�;�1h��˪G�O!fy�-Tn?�c�&�&��c����6��r��)_�hSK�s����Aw�䃣_�xS���x�˵B��k6�3wyRHn�^��p����^�����u�'��5�K3����+��;k:S�;?nV�X�fB�����S��90�Ԓw�@17�t���^�fg�{D�n40'����WVjv�BFh(:#���$�A�:��ظpwC'2cu��̚沉����&q>�`�JAj¤��F
������ �9�	n�$v��g"m��=+ޏm�+s�������+��OE�W�j��0g�WQz,*��b�ϕN��
�ʰI�
w���G����gffĭ�h��^�9%#��)���J�=�f�N��6C��d���?�����E�;̐+�� ���4�8	��3�C8Ҳ;����F|���3[(ޟ\������g������c��^���.����\�=��[�rov���(�����Au)��6�d�Z��N)� 7MCl��� S0%�Ve,���:�Y��sa��3��L���{&��ߌ��{v 1q��ʼ�fܴ�]A��4>ԉB��r������	�	��Α��>�k�6��f�&���^��:���V�_��Yd���h�v��N�~�6�da+�j��.o�����E��+v���k��Si�8�r�К�P#�������r���+�Y�g_���[���Q;ntJ�g�)?�gǵ�Y�.v��c}�C|��ɕ /Z$�Ci��lz@A!c�����{՞ns�r%T1��״��pW36��<�g\IҼ3u���t̃�t�����L]ڰQ2�ݘe!v�\s`k)���(9l�Z6Y��(?ں����iZ�����Z�7�Gd�}�ж���JM{�y�'�D���"��=�\��f�`[k����{��W�Y�<U�D�~�������z6,����n3��� A�[؅<7�+�ܕ��=[�
��<�ʥ���y�*���i�Eȗ�zng���g�#l�pz�2�1:Q�$aX'Κp�k���=±�΢ҍj���U�P�� +?,w�!�ɋZ_�����N�����	�.���n�W����4�����2���>��\����=Wx��FQѹ��hv� �<�6+I�a'U���,��g�sav"���{F\��b?�*��{����[�GY�e��pw�����1���n��N�տj�-jƂ�:���-1�1E�G	�ÁQ���e����ʆ�w/�-��0�q���V���:wa��g�|����y����-̰r���t���`؅FXy�3�����sЧ��[�;��X��Hk\�c��>�<=ۭ-uA�1�I�J�x5�a!U���՛{^�Y�e�3I=�w*��.��i�?λ�Af/QY�7�%3~���yv5I�[W\G�$s����4�~�RWUH��0�
WCZ����G�������̆[Ƨ���	�[i�-n�GxD�n�*��<u�H�5�\�;�\	�{�z�O-6Em��j8��i��ꍍ��7Ű���͐�����E".�Ń�:TdCqdy�����9�2,����'_uǿ�TT�H.����_�+����}��Ӭ��_B�յ��4"Ʋ���"gB],1���x�'����)� ��u���)͹�Dϓ�5Ӭ\]�KO����%�YM[�3�	��)G��:J���p��L:��%�c���Q5"�9w<�R7A����xn٢����"��+Ո���5f���@�8B(b�2���p����6�o4���\���@̪��/���<����f���w&����a+}�h�ڔ�m_r�I��t�%��3hG�d�Z��u�p�˩�2��#��ۻK K�>�qK;�D��&�i#$�E����V߭�'��*��*�"-���h��t�A$�pC>eU����p��Ap*�{)����2W���*q���3ޟF7[?�O	�C]\j��t=��6����ͫ�����X^k*Ə���,��\'c���B��M|��ZJ���`as���'\�nwvb�F��/<e��A:��cU@�2��=/�g�x��~2��8�ֱ:a}J8��g�$��)�����m��,V
��2}�'���b��@=��om}Z��έF��F156�[-'�������}2h\��?١�O�00���g7���!�5����u��b��)�+�$C��c������ȓ�� �ZD�
�#�g����Fr/��u���(T�:����s�p�[����ëa,����E�q�7�$0j�p��H����
�Ȼ��OZ/�v�*W�^��5�[�B���	�6���"z��cR�1��XB������j��l�<�� k�/l|�t#��W�͎�,nV�y*�
4�Xlۢ�$��U�m��}MC����_\Ot��������>��g�`���b����_ʋ�\�ܸ�ǯ?��Hx�Ny?dڞ��Wu�|�Pc%��F��;f��.E��ty'�Ɔ����|D�M:�㔗�_�e����$�I��+���,���̾s�p���e�k�$:|LT�C�K�)��������o��.�| �flՄ�29o7��Il�����s�Ћ�d���zM��R���?k9�'ö͘�$����M�5i����[�����'�?�@}��m�w���K�lbkŹ�w�l.�'�A�W�?�S���>�?�2���0^<���%E:O�뭁'�Q\%�%��j���x"�R{�a��w)��l�.�3=ny_��H��	\�Sz�����7��Ч˳��\���,��Tm��f,���V��M2g�p2[�'�������
�N���Ob�/��C�/����k�3����>xŖ�3���(����e�����6�3{4J�/��h�iDy_��ʈ���W5��9�X���D��7��2_��h��@;�hh�9�*	`E��@�X�|�H֣��+M���1n0��͹�H�|�E(1���v�����n~��D�m��Ʊ�4�;�y�>Kt1N�n����=+��Ý�e%Ohбw�vk�Ѐ7�b�b�(�򂶵RYScH�Ϯ��	Q�p��#�zV|ZVܼ�;Z�`�+*�F�ɩ|�%Xd��;L�����ӵ(�! �vM}X���\��X��yJ�����u8���6-_��x��s���4�D����[��1'����hc��%�ធ���&�3d�sx�1�W̧�) Q~F�V���m�7����ϕ�_�d���_���z3N����v����q�s�-�V���d���g�+jڋ"ĕ���=h%� ��B�A����G��������HG��v�5yq�-7���B��r���9�I����)j�l&����	ξ�P/���C΁�sXP��ŖI��E��9��2�%'��`v7H_V�{ǅ�w�L�*�Ɣ�>�t�<K��g�uq��*nr8"}�~�{+\es12��T�I�8�����8���qI�Ut��#+�5�y�wv��k��0�O.�n���V��l�//.e�r�������r�$�Ɨ{�!��h��.{�G���r��?�]ޣ��9[�Ns�[�_����);�:,��j�4��T��~twy��ΐ?�a�r�t|t*��{<ud ���t���]�n����E Ua�_1	�C)ف�b��]�Y���n��XMw{��å��\��J�~����$S��eEf���9�S�ɗ�M���/�>�I^)#gI���=)p�]DRyV���sW�ĩ�q�IasZ���u.�Z��a��X���Ј���c|�b�O��K7*性��e�Ҿ,k�0䚥�|A�Ҙˍ�}�KU�t��m���C�KЭ)I�'�5W�}�s���9 ���=���[!`�7fA	����*�`l2��T-~<F�_Fh0���%#)�Ά�Å16v��w�������D�Ify�C~�1�JxR��I$T��	���<3zv�G��������ox,��{pPna����5p�υ���ur���AXK^ل4V8@��79�B�X�&^���_PV�ۥ�9;��&�Kc�'������S��Y��\����jc�*I0+3V��g�j��K�g��]8!B�E�	p�7�m��<Ί~zlɾ�5-�d	����O�YvM�>�f����靆�Ew��[ޭvܲ�-WbouZޕ�q���%� nWҬѽWW�������,I��w�Kw 9��=��[��2'�xbdϑ�������* ��� ����������U�c��IeKO�|BN <�4���q����L\��T����2�~����^8�q�.RV[�<���]`!E=� �N�_�$�[���,������	<���ht/`'���e������R[�1�-��o�"*�N�k��+���ٓp�D��M��ɕ�#�g����vY�VW�D�����Y���M�B�$��W����>w�a�(���T/@`���B�84gزeTΑ�K-��.ǃ=
��c�pT���vt\1���5�g]�������G\�� �}7(7���̅	�n���"�9��/��ik�/&!`Ӻ,���,v�����8ƍ�q�>C�'��Z��P�����J	�zG�?ˁ"�Ν�#��9-�-��R+�a.G�}3��2u8��9�b�_	[�p�8�H��-�[�C^���nX3+��9Q�O�o1G=w�J��[�F i����~���PB����8��F5�V~�:�b�t��Y���e��*+������Љ�Y���=^����`V�O	��+��X���
+�]$l�d�������� �� ���Ȝw;�pI�u�7U7�Hw��{�?�Q�ʬ[���/ex�����q�� W�vؽ��&<z�o���ۚv�[=�K]�]�@���Eӽ�_^�<��>T<w\b�@6HÍ/�I�V�F���KGW��6~�����hi�*	\��u���uM���Ž�;��4_�Km�XMz|�)[�[nN{���O���i+�/z^"a��~d��L���#ٺ�iC�}o�<�-�W�N��;8�}U�ÅS�����7�3(1�z#� -�����p$W��.�����H�AK��Mn�`��bO�4�1��ٿ�5������d������p�4s���Ɖ5��c��X{�Fi�cc{�:�B�{�fc���[ �p�,ꅘ�G��L�W��	~k7��|ςڿ�5~��~i��D��������Q��2q���mA�Y�Wl���ӳ]}���(�)���z���_W�p�IbJ���U���U�}q�U0/�n �K��O�/�e������zl6�n`	N �iE�03�@r.�Pd�+�b��í������e�5}�ajby��z��!�t|u�	0�+\�ѧ�~u��eV��i�3��ox��(=��V�o��Vצv�f�㯱Ʊ1���6qS���k�h�� �+\nmq�r3���/�d`������[���ڱ���B$���~��k�Bx��
Z��źZu�W3�r���σ�m?��Pj�=[;۝nv]{>[e����f;I��V��4b2g�U�`M���&�ľ[Dk�����d$�M-������A �\�����ѷe��证j$���^��gU�&� !�&���Dk�@��}D��ٞ�UبF��!�Ƨ����m��	�sL[��H��I��W��Y�����*EA�X*5�a��{��u�;aϋ3�|ˮ�&|��r��HD
�k�fp1M����4�,W泛��&)�Z��;nEn�,�­����	̺�I�6&S��	�gA�D+5������rL�mv��5�|Y�_{\��A�s���^�gG��h��}P�]�W8���Ջ�5�*��-��'���.��Z���s �S����Stt7�;A$#��&�u�G���[��}HT���(�!L�e/Z����H�_��{���%ԇ5N���W�IyI��)Z���O��J�b��>��������R�K������\Hn���z���G�}E�ihf	��	ש��="�p�Bu��B��]�pX]�y8v�/�A�@����X'�M^:Z�r��*f�T5�@f4��!�y����d(�LĢ`��a�k��b�+��%�+Q\DfT�e>.{?͂�
0ک��J���x����8�ؚ��3*cć[c��?�A*)�����a�������6���y�A����zE<i��U70!��I���!4�Hw��4��ݣ�;���;AGN�ֶ��M�ogg���X%955����g�(�x���0��q��冱8X�z��f��{r�>_��Ķ�1��y�m�`a�9��lH�8D[ϓ/mh{>�$�����ً���Lq^��ǒ�t��:��.�3�d�Ę?�K�YU����ԄҮ��'K�'�����-�5�D�}
�t�pC�'M�0@�"ڟ�U@\$~EĬυ��&W�b�����Zwor�_����a.{,�z���zmXJ��,��x�˂��cr{,�()��I����}��'���[
r�OCK?Re�~���w�N��-s�X�&�8z�h�~Gơt}x?�v�wYg=�z�u�"2���%;}D��l���~2[Re�`߷�RjWjk�8�FiP�+N��5i8P���]]t<%��z�&�3�P�]�4����׋=H�֘�hW�E�c�p�/��ċ��˼��%�+;��Rlۢ��CD6�T4�2XE��o����t'��bg�h�Xl����<��J:���o�S�CI�όJ�+=V�.���Bw�b�I,O�gr���,끫ID`۟��@)�걟͹��1�[��k�u�ہq��|u��|���A�A��W�L��T<��ٟY$�B�7�ᔔwDVzuYxqx�A���dalln ���d	�'����^�-j���޺ݤL��{Pb@n\��6�Q��+e*TI�Ӓ�H/�_)����Z��p�O�����?����܈�V���b7ĵtcW�Y��6�9�Oh�2=h�u�F�a,���I�K�cZ�c5����s�I����XD�5�bHٟK���	Q�b��PA�%lXY�tg��c�S~}� ES ���#Wd	S�if�ķ����gY��I��\�
}2S�R,������P"���F�(3����m=���"���ʋ����Vg�~�{�����j��ô��?����h�"%�������Ę#TqK3�K�C��B���q�so����p����v��,��Ĭ����?+hBK����>�Y(=V��MB0��g[��r�Z�P���8�L{��|�+�'��;�98���ߣ]�3 :,��7����2��*�ڍT�	F$.J��mJ5���gJ��zpaU�zs՜��\� w��M�֥���Y���kL%]Ms�?{/t�7�Z4�K%)/��,!��|B��~�y��p�)�F+%�6z�r$��y�X�ȫ�osd��"�l���7f�V+N<&����q�q>!������*��8���1-`Kx��y�&�{�)|�g�J��-Ye�[Q�L��;K��.=�����G��$�3������
�hV��n��-������+ss��-m�o�a4����v&F<ݘ��vۍ�ia{�U)��g�	,�>D��f�
e��gPdVSp6��_���K�� �����Jf���7��� ��6N:�Pe{j�
�/�B�>��p���~�KZw4''��R%����\)�W4'~���Z�.�}���E@�_����a�=��A�k�>c[�4-n��S�؋X���{�x���a��4��"�7g8
�L��ؐ M��B[��VB��#�^��b�5�s7\�U�c��B5gDh�\2l�V��<�U�p��7��� _����*����-�m�Fs31R��5?�:`_��.Г6!#�@������u��P��xNω��$�ʸ(�E
��г���eɓ!C�"q��z�V��q���A�F�����	����?��ݒZrx3fV�s� ����5R y�@�������x,�&����Q����	5���#�~�9Ot��2��_��ܘ&��_�YG���"}�'�k������_� ���19oOv��YX4/�98
�B��g���b5fϾ���:~��9r �qB����'1�]H��b�����XLL.�9.Ķ��g:z�����L��R�}������7��4~�h�Qi���[:+�#;l
�|��q�������2}���W�c*�~Fd��5X����N�#�B,��W���~��/�����P�.��<׊�a��;XeM��6��� ���XlW0 Ӫ6��U :5����gV#h4G�!R���lc$`aʾ ���ί�u?���K%Y'$���>S �	נ䳺`ᣞڎ�`-�w;�A��v ����F@H��f?='��׆�^�sꏕF ��p�e��N��]����lWИ6Yʤ��
�@<*��ῐ���޵O:�~WR!i�1Uv��WG������ŉ�z$�n����Bj����o����!����ڔ?\�ߴ�] c�2��O�P_䌏{����ϟ]��0���W�7�����I���څ*����!�!c]���7zhl�j���	��R�A*��~m���^*�a�+��>�ja(���X��NX>�N�xb��aA�`t�.bsz�:�"����^{��;vZM_1�Ç�$�vL�� )!�yc5}��W:��c�JM�k�����VV���27�t��,[I l�sr���q3�Ek�f\���Y�?�@"�2�T$�Hbig��=���.�L9�}@-LLe�DZ��^�#��O������Ո�w��v��2� �~�:B�-3�^���!�ԕ-���`3��C�N��"tAg�A�EVY�B��ҝy2~���\�K��㱗,�0{�}���iʻ���;���2b1���G�ҿ�ʹ�8�?H�r�GM��g���	�lP�  ��/�/z��2e�^��3�$gj�K�8-�N��2.����ђ�! �(��y��&ǞN�{��7�ק>���ݍњ��[�æ]|�_�tA�����A#]Ɛ[*w=,:^~H�G�A�gr����a*�űG�mZ�g~\��^��\�H,��4~e�w���rqȺ�Ե�ޱ��R�F�`��ɦ��-`�㭅����3�t��|��}B-t���G�I7p��
Vm9V��iaI��?� ͋���g��_5�����cn�1u?�����ňk��E���q���;@�e<S�_��O�Hh�U�ڔy:m�@/V�ߖ]�O����RD탣n$�J�Ԉ�u�J�YW	���=��6��Q��̈���e���\��=P��[c19���*��z҂� �:�m�ҧ�v, ���*�2�q]@:�va�F�K
��E|V��~-��F��i�ࡪ�x0R��ߊD�Ws�`�F�'T��|���������9�r��_�T�~����q,Q,r9G�����w��I>�G6���K�wGD2X].��ĳY����Xۜ���f�z��K��������!(?|S��x����oTR�"��~�,�߆�Y�{_�l��07��CQ֜�ќ3v[n8⫆d)W��1�m~n��;�������X�]@��8���m�{���x
!�|Z7zHsQe����o�14勃T�����F+Xح�v��>����Ԥ�"���c�i\�-�����y���ZIM�
�������_�UEG��	���Dڥc����3W��F Q�)nS�G�/���e"��m�tj�c`ﾮ-�~��%1�m
��o���r25�'y��9�~�S��\�$�KE� Rlc|��{S�Ŏ1�lًjĤ��X�ъ���N���1�]J8C����G)�=����ym���Q�0+��lϧ�+����9�Ɂ"Z=Y��8QpLR%����p����6�|��s��Y�������kr��L�Lrr+G߰��߽CB�2�W�/����_?����o����^�I0L)Zcuw�X|�?U����x�0j!-ꤐ��BOc����\~8��h)����~�_��&h;�b2�F^">�^&�,3XW�����,�+ݳ���ʺJ)�'����e�{z����C����P���t/K���Q��������~�:��
U寪��^E��c��4�l�P�;Xgs�����ְ�\�&?/�t��I`�t;>f���s4�cz3Br%wЬ������QV2c�$T�$�����NםCKM��x��ȫ�Mޫn����Rm���n�<�:X�@���/�L���r���Dkd\�hT�FB�p����"s�6 Z����}3Y��R��j�<Qـ�������ρxڨy�W�C�>+�E(l�\-��"�D"��k�Ir/�+E��}�	"3��M_�7P�ݔ1�	��	&Cz�߾$P��^�62z���xȵ��/D ͧo�d}�d�4�uyV>z&v�%3��:!��t�l͔ä���Td�sR)G�l[W���bF]:��O���Ў�L� 0Q��2�6ti���D �q�ُ.�������(�����Ŷ�XZ�L��aX�z�|AV㩲�4w�q�@��ƭ�l��¥}'��~��i���D'���A֟�i>��l��<��U��[��cK� �,�1؉;O��r���+�����0!�lOƇ���F�R���d�k�T?���jIEK���OC�a8�H�
6S���]�b(x[-Hx���Zl9�������D��t����-����ZjQ5͏�U�zjuOUr\i��1�H����U��/	��	u��ʿ��݅#��f{�J��dY����J ~qËuFT�.f4#K����C<t|,�� ������7� �h|��7|�q5>��%~��IX��j��e3��6#��0��+�2�`)��i���l��i���GL�Z��cV7�~.�!k\�B�X�4�����S�4����
D]�"Zfm������zڲ�4s?��L��9R*��=\+�{o�͍��NԈp���Á����4�rk:@�/�m�1+�8@Z�J���%:]��m��u%ݹ:�f�J���P,�g��w�����?��/8��
$��/�ВC*s�vI}ޯr��m)���J��w�a�e}.��=�?���(ܗL�4�� VZ���y�+oLH �76� y�jqzv6�?�e�y���"��ӂ4��ܭ��uɛeR�����ʅ�c�}T#{پ���'� Ӟ���H�)�T�}��B8��)�e�B�5�v��/�U48ca�6�ue����l��_N����F�n9d�t�K \�-8�:��lܤ��!c�G���p#�Un9���&�A
����j=�������� ���9�F�$����g�б)�}�]���(��7�m�^�p3ت����:�Q����3��Ǭ�r	8̒�J��dpfSV�ҲJv����/f�3^Y�rq2� 9�)��εÁj��ͨF�X�D�xg�x�^Ѣ!*5P���&��f�8A��JSȟc���h��y�*v~E+y�o�Nz�����z����QVg*�7��]�Ku��
��	giii�k��iv��7_"d�9Kq�+��Q<Ԟ�}]
Y'm`�S�X�llLj?&��lq!�%ߡv�F�ū��7�6����66��p�z�Wd�⺸�_�c�2F�61���C�����\��ѯ1pCg���q��]Lx�b�׊��y�RDR/qa��NI��]H# PV^k�7���Bb��,���t�����2Q�|}��Q�����5&���$j��R��4�x�h���.�^�"ۙ����DJ�?K��&>������7�,ٓ�h\Q9��"��b�&�i���|���)��<*esL?b��t�����M��t7�س�D]R"%^$�����u$[泐1w9���YcJJJZ��X�.��n���C�S*
J���᫩��I�u�U�����Wڢ;�����DX/�Fk�rat��n�g�z/��{�~�t�*>��NFf�"�.�����B�\�jZ�1l�#냳oT�_t��ĥ��j?� �vM^_���`�u�	E�H��n���u�i�=���X�0��E��9k�}���i�h�*?�3�#������s�L��x�N��U�<�>C(��U�eV�e3X�[a��O�b�Ⱥ��l��}h�q���l�����D��W�S
T���GվsS��]��+Qn��/�<�p�5�Y=�g
E��sM� ���vm�h0�)Zs�t\N��5�@��K_���kV��_�w{����X�}ץc���7V��cV�b7��2?���,����Wc(��*6�j��^5���C���6`�[����=`� |�	��z�D�}c�6�����ٖTLt�����]��<��Cm�Ƚ��ݟ�,��RL��b�doTc�C�i� J����b�(G(_-�p)���͑t#A�ߓ�W���s�Ϲ5�6�޺�E�����dm|{��E�U�.+��&4�3�\ �f�	����Ⱥ"O�P�%�:D��,u_����E��e�|��2Y�
]G)�7#�H�+�>k�= B�-�����gU��շ�BFm��kױ!`af�wsy�����9�poL(��K2��lݪ�c��M� I���؛Sꥇ���$��
�}��q��움]�b5�,Vd��O��)||%###^$w��;*v��cT=�(�4>P��hP�P�m[��h��Jv�>g����[��tq�Zi&���c�W-�iR���
�$ҽÖ��]�b�
�
�,������5(>OMAD��-�ck��qt�Z<��f��������.��O��By��8�A"�6�:)�?��w�>���wz��z�O������~"�d�J�u.��������'թ�n��谏`�qJw3���_�A��I�>�~�mBCH�ɽYEP�,Tr���]ѐI��>��7�ma��%�����<�d�z�_!lT��Sseh��͒��,l�h66>q�$V�f[�� o�nGm/qQ������]�tw�����
?�V�<��� ɕ����@/c^�q������P��t���z�k6W��9�?�oovC�CGϐ�Y�7�(�z�hL�W�h��&qy���=����=����>�6�,��_?Md���#Z!�S!����5�Nf˟�G��q�Ad�x�
>|�>���@/��o��/v��6��I��^��m�-��ԈVm�	q;Sn�o�e���K���d���4�X�~��#���)���]��#� �ˎ�8�Rko�9�W	�b���i�\cΓ����KY��~�N�D���c3��H���41k��y��P��NZ�r���!��m&×N�2��J����Dm����B�m)1�o/����3�^[��Ϩ�?$��?w��m̕@j��΂s�f��{k�U��n�M��y٪��X^�F,��'̸�0E�AW�~[�˱�LdM}�����5b�O6z �AJ7�V<nVS��5���K���������n���w��M~�|�o�˳&u������ժFX�@v*� �|δ2��Pwl@��X��y}�j�(�_F����+�$�
)���P��E���� �)د	^f��(d�zp���a"sJZ�;H@������%q� ^��~T�̴k��)�t+�uI��5A����smΨx=�Rl�(D�� :�1jU䡴��0I�
ko���Zu�<"�L%?xV9�z���7��B;�܋�P'I��جZ�����UZC�uEͨr�����Χ6���mkc���^A���c���6�sRo�=��mE^�HT�4\���͠@�G�?�ޢ���oV3p�����L�&dKK��aI��P��R���Y\d�Y+�W��D��LF��hy�`� {W����wq��1�%@sp`��黛�2��[��UwSpu2�s��.��/�9�,)yy��S�m���W���/��.�SZ)%��~P,�[G����d�5���!�ߍ����?�V+�_^�i'��y��Y�6��?�ߥJ �+�� �3�Yorp�!Ⴢb`��4纾�e�*/%K�kҏվ���ZӽY���O"�"o�F�9��B
�;��_Wԛ-�)�?���$RZ�.�n�4򷌌�,'w��B�E�/���/�B8��bͨO��H����$���(#>oln��Xw7�2�A�{�){�����5�2���gCnN��K������ ��� �3��h�u�*�Bdy̟�1�&����8[2"���`�稦����|b�f�²�ⶤj��i��j�ÙN��_:<f)��|PPЁ��L?i�׻�w�Dg(��fި�Y�?xT&��*x����fi��2�^?�
u�����0�_A�F]�q8��#E(lg)�����v��Ry��M�g���Ǔ��c���H���UPQ�B�u��0��ݎ ������dV)��;eQ^�S)|�g���[&Fk��u��us�ß��8O��b��D�]޽sx���o�Ҙ���j���2��/�-�ٿ����s$<�H����i�!����Ki�\ 
��}i�Ł%�@���Ë$�ۯ�����O7��L��*zw�O����ס��'q4D���$1ā����S�uj��s9F���Q?�g����+��}=Z�[MA*��WN$��0�Bm8�ex��P���W��ۖ^.0����<���X��g�Մ{SƆ�n�Z)�=a�c���Y������R���lh۠�:���[�ڃ�C*�i�!a�Fłr]�A%���R��oVX��x��/�>Y#/��~0�4�H_C���7�:����ٝ�$d!��..ˑ؛䁥��=<{��]��׫a��-�����>�o6s�5ro㬟�G��T�R���*K��G
J�h�;1Đ������"l���9�V������F�B�� Z-vG^������yI���7�GZ�Mx�7;���q
��I�+�`�P,L��J�4f(�?���b&���;.3���Ѯ��W��@φ����pg'�!}��m��ߍf`ApЕR\[X���mӝ���̈́_�n��@*���j�T��DK�!wk[�3:`���Jʮe�N${�p{dmg�q!�q��m�șo�!0J(�vx)3���4������[��l
.顨6���.1!�7I�V��R��8�9�_��M_jjͷ��?��3����{oѓH-z���#A���E�DD���^G�ޢ������{}g�������>g���>{��hM}�nY�0酜�� ��Q��������eK����6��G���	���K
���Q��#���Ir�'�7��?+��`C��c*�}���ԟxz� v4g�KE�&���k��q���UW��q�{���_�ld���w�%2�p�S�>��{X�xA:Mڛ���2V\�]�ꖕ�{0	<1y��o�yz������	Q���6F��r}����u�8Ib���b��م�����9�Y��0_>�鿪��*h}��lh��
v՝���{�a�حƃ�J��8lsL� �A�W�H�8�LM(�F���$�����J�`MQhN*�����ɉkso��RS_/��9ѹ+w���5�����K񼽪�C���_��_��[�P�e'�e�餳�f�����LD{�\o������Ǉ����V3��Z�H�o�>��ײQ!ڶA)<` �ŏ��ɶ��e.�����ן���D���IvK֋��p�ɑ�x)A�/�Zin���m�'ci2����S<��ñ���z��MS>�#q���#ҝEz�p��[���y�r�`�"/dL�8�N���,����n/�t�ղc�/K��zP�����o%��:��x�j�%؍� �V�̠a"��;��K]T7�Aᦱ�;b������P������dY'-L�w�@[:&�����&%��+�V�fZ�'�?�J�z��ٳrM��[���){�Lju|/����K�3\���Nd����R��|�1
��a"�z׀�J ��Ճs"K`m�2���G}���_�䴡ɔX7�*����������������h\����qR �)�/�p�|;r�o��tص�e�ӱɃ����֛�}S���JFi����w�����<?M���-�X�H&]�b棉�.��͐�>���Z.�)�VU�z�N����$�MA��bykC�!���@xN!��E���f�9���4�҂z�rJK����1������;H�e|��&�/�E�ȏ��:��ೳO�<i��ߨ����ӣ<::z]C�C�TPP�<ۥ/.)Y�9;;yw{u�,�E�,���J���#x9R�UY�R�&A�����&<{Ϧ��~G�4�:��J(��ۡi]����0�_Z������|�_��;W�6-���x,�8�8�T����w١׫m915�o2��5o(��F!'%�˼4�A��9�h�q�3^��)횭pt�턲�ؘ�D�����ls��QNlu���!��$D ��k������ ���6ʒ...����[��=N--�Q*3y�� ^���Da!���(ZR�y~͉z�?\@(~���^�fg'��{/TBb�	+�B�*Vf�p?4�ef`�w� ����n�g�ms��g=J�sx|�GDJ����ʿ�ޚ��-���8���%3[�ɯ종�����{$%$F����y���x����y�I��B5�_y/�F����`pBb������~O��^�/t��+�u�10D��奲��i�����^	�9�3$����hu8XW��S��j��X_s6E󇗻w�F�G���kdX���"'N&7�(�׸�n#�$>s�� ,;���|;@c
'٢����`s8s-��gr�3���^N�Bܾ���~L����k�:Ȼ�k�:C�*�Tɩ�6M�}�<ݍ�	�9����11�h���6�|��SMъ3.RM,�$,8rd�F]��6:@`q�b�����n)�*�8�6<�+Y�7u�7u��я�U���g}䎈�.Dsd�O7e��/ ��3����4��mz�m����߸�^������{ ��Zh�|K�u(ޗ˔�J�� E�$)�(��ǵ�Pg���ǿ4�����n��NHBW�=,��k�����Q��T~g����r5Vr#uKR��3?"N�ʶ+j�氧ɨ1*!>���x*>U��jgdW�}�����J�r}�,ٚaV#"j�{Je>{~<;1�jA��H�b.�<Uf�Fn`b�(���\);��2���6��K^K+�y�De4ۏ;V�|���8���9F�4���ϣ�	ƧD�>�*}��S+]3����~mu���ĕP��\�����󾤤���­NmzBB*���F�b�݁�ZZZ��E�s���?�v�B�b����7����yF�B��T����D�M^�	t)
�t�E�.
˰��+"nϾb�2����`�7��K�;S�!X�}����0\���u�{aZg�{tɸi���]�x�}c�wXi�����@c��ø�'C��*󋺃/ͺ�����5x{�	`�H�<id���7�pm���KeTB6
�#֡�6��;l�b���[��H�Jy����&��.���š��''W���> ��k���#~�q.�=̬�U�Q���[m�9��=��'~Y���[��k��D��*�^д�qՊ����e��
Z�3xun�2]i��������S�X��|�w�_��o	��a\�DX�X�%$�n��M�*M��.�ɷ��V���ř�ô.L"�F�	i����x�Z�1���V�m��떇�~r�
O�-I��!&��w�^��={g��=�������#��f���QVW~iB[�;����V-�kg�:靿UL%���AV<�P�_����rs[�a��G)�~����V ��mp�Lq
��ފ��v����N�w��K�t����U.���u~�wH����dSq����,5[=W�hM	�[�������mO � �Q_R�_�@�gs�w]��ԃf#�sw����J������f/15<�?�.&�uc}y�.�� ��NqI~��0�P�c����ٞ��2�S�G� h�AD̊�N�;`������mvC�$������g�˔����|L���D8w������;��b�diGH�N����*�\��K,ܴo:H�ј�^;3���6h��K�g
�C?��u�֨`cUz�jH/��W�oV��+q�A��*�s�tp�TQL#j2�D���̺VfD�B��k�<������W
 ~W�����.1I�T|���F<z�yMb���	�y~ն�C'��뫊�����s/���S����IB�]0�;[8q<��q�FGE��-� �ڽ��
�HL3酩aS]�Y�WߟvA~�6[QZ0�-EO�ƍ��s�c�T�"����s�uT�����)<��'BXm��6����f83.�	�Em`�j�h6�3�c�˭�����_F��/�z���vgy#�	˳ù�_�{�B��/����Y.ꤟe=�	28�=��貓��`�T� ��~��&JT˨`3H�}u�;��η��Q�E��@�zv>�4

S�NK~��Ws`�b���1��ҹ;(���#г�8�$�|�e�0y����&�*�|�'��G4�q��:�Vi=����I.7���/�qŶ	ևZib&����OV<A<w��)t��Y��[_���FD���yH8x}�4BDR�S";P�"n��;���G��X�!��(�:�3͕�(��o���&O'4`O� �;�^s8����uv$l�:�Ď��D�gy�v�����"رԅ�Y�W�i�`���1�����B��|�͟��|��FU�kjz'�^c]T����w�\���?�:�||����k\e
��}�(����T��뇽c�7V�վxϣUU�m�L�x���`Lpv���U_q 7�6b��W�����_<��	)��[�u�����п�-�������{1O��A^�����O�Ž=u��#��?��Q�Q��R�x&ɄZ:��+�Lsh��L�\Z�'��7���Ik|�U���)ڣ�ذ���f��$�^��i21g��Z'�#��������׀���>W�s�7km�A��ѡ�8R�O�D�o7�bv>bk&=A�|I��"�<�m �u&0�랡�o��nu����:�f�KZ��xEX���{��
Q��a�m����C�-�t;�e=EV��B��/Q�ᔐ��8^��g��Sşp^�މ��t�����R�bO�t�ssv��!	{�Z'Y����06jc�q;��.��Aeo����w�d��k���.�:�[�Cm�3�Q	}����-m2ch�n��߶��%�\��?F&~��L>|\�����f��[����3�+"�����(Z��_��Ŏ�	�=M1b�\�/^�(�u����R�2�YvnK�|+�g�T��n�B$��x��H&g����h% h`��D��ﶷNN,�"���`?-��N�b���y-�t�.,��s��}��H`�%����&��ٮ�3��?e�_��͒B< �}7�����; �g&qN	�b�G0��=m	��Y�������q֨�~ei�7bIE9k���'k�F�������P➳���Ew��HD��j&Kxx� ��2ݚ�8�/{��5#A�߰�y+]���y���I��3�}��/�l��F�� �$D�O~���W���J��%�&�?H��Ox���I7��,��+NɿJ� �#Kd�����D�����*j����d��rE��A��	�Z/�}��H0Z#P��3,>��7��DK����_r��,���9�d�L�p��X]_�J�i�ãP<�q\��s�~��S�m)\��Yij:�}rIPyDр�f�����S����{�2�S�$�NZ�Qڡg@@�"/�Ct]�d��t�V5�Gڜ)�i��Հ� Zw��n�z�����q*=3.P-��\���`��W=���,o}�`�6���������"*�_s'�t�2"�y:4�b6r�ik��Ͱ��S!�Ѐ��	�ah屵���Q�cQ���4���]G���!��	�\�%�Q���p�O�J��?/�'�-S�vuay9�*��6<҇�n���!	�d�������9w�&�wJO|Y�$�bw�a�(�y��H-�����|bp7s����@����*X���R{������Y~y6>zĚ Vǳ����F������Y�ɿ� =�(���Qg\�m��Q!+�xDb5v���x��^ ��J��&���j �jqK�fSƿ��yC3(�؁8�Jz6�̕et�_s;���"�7!�uT��C�!6�~�{1��j�H1�����[��;`탬7t?~�>�z8�aq�{u�7� �o�����Õ�f!T�Q��_�R$�<�*�u�z�W����/�N���)��z������Y��&���M��X��3�P�">��0e]�+���00�����M������6/ND�����B%��h��I�d��`��µw�C����s9��X5�B�Z����~7���?����6.`����_��"�1���n�6~�����\�Ĩ�&$�?�U�M����Nj��CAf)�%��r�z{��0��%��ׄt�2���I3.,,EJe56�P��At-��F��4�&gg<����Ʒ���²�EΧ�I��<� �(h�	��$k�sB�)�=$~#���0���7�9�/�q,+�c9��ʹ�U�.��/��E�S��0�P4wa���n��mFU�m�b�>9n�ց���ި�@a�����(�P�X�l9��JQ�B�2WJ&�������L�H�>�ϐ��]F-�9�{�ɾVR�?:>�w���s� ���r!�|:�aS����d��s�rR���S��I�Q_�L�yc�)M��i��n�6f#iqȘ��ܙ�bO_���2�����ȟy�8��V������s��fۤ^�|��Q_����*3�
۳��8���6#�Gl�Q��t�����ŧʋ�:�:�@\(��RS_�s�%+S0�+Z�B-�Z-�d�b���\#eggg%�o�[O�ߖ��&�LG��$A�G����P䯞mb���23GJ�*K�ﶟ2�l7���	qq7r�Q�[��mMz�~ �?�J���W[�"�X1rL��6%㰔V�n�����c3�=!V�����t�(��.�T�P����uض,�D��6�a,H2� �������vG7t�ƒ�M���ݙ���ȨH�5�v	ʝ0���zT7D�a�K��L�SpGQ>�D�eJ������ ��(�p��1e�9�>��b�N�N�z�N������I!�3c�/zb�<������V��VPٞ2�������b�����5�k����@d_<���N��^GlƿvHRB���#E�Nr��:E	�$�ϟsw�iDO�kp�A�L��±�'W敮����֘�=��;���jHNN-�d���D.�j<e`B�8��ۡ<g����>�/���V�a�q�
��}����FF��O���A�^T��{��Xg�'��#Z�}+��|E�m7�ݧVkE(�YG�2S���'7�SC�.S��j%��^�u�[��<��;MJ��A��rr["�Q�u&	 ��G�;��|�;'���s��Ѥ�E��D�����Y��؏�w��O��o����g�G�֢m�D����W(x=���o�e�JӊǙ�������A+}_s�4G�ʁ��D��OH�JɋBŐ����M�x3{��*��}ʇ�b]36�Y�D�C稼OTm�-\]u�
9J1ҞK�����=��l�����ޟk��O��G�}b21�#d��Ɵ�R����KO�o
������Q�m-�����M9/��l�|:P��ނ��݃?<��q�VB�RPT|��>���~۟u <�"����ayE�n��2�G�~�7U�^b��p�s����xr�E�sw8	�����?��ԉ���_F1�����T^ؙNT����^���:�j�p�l*A��o���;pK��("�ݍ�w��i?x3��F4brfU���0�1�ƈ�o�ؒ�� �*Ҭ�b*��Rp�03{�k0={z���%WA󆳺��톂��L�����Ǭ�h�i�Cj�H�M�fǩ��$�t�l�lϐ��ypu�=��d$�ӱ������5�x��Z�4���8���4���AZ��dlޯ�%���Վ%{��&R?��U��o���x�B�)�@(8~T��
����'+}�P��� �AVzZ(�,���_�A!Yx*A��]��d%̹SvOP�[��A�x��k�O�)���@�pLL���LS�u���W�6��im���������G��C &��9���YE}/]�o.$BAj4E�y�Q	�6�2U7-�a�sk�2R��P��fIYV���EW ����wzQЛ�����6����i�䯏��&�D��֩'d��
ˣ�F�P�#W�Zɦ���'Ϗ��y��rG�@0^"RR�XN]ug;����-�.:E��'x6��Bg���{P	����V�y���=���]�k�~�i���Aibrk'��1:n&ߧ��YS�):ByYg�҇�?[=l�A��"�5���!0k
�{�����o��H�[qiq������ɷɩBڃ!������.�.���R�u�X���
�:�f�ĢQl
�� ��Q:��\��[	H�Z�����}	��趤|�P<!�/R+$G�czT�j�>JIύ�B����@�dI�.�ܦ�&���xkC1rw߽]-���]�4Aġ܊��|Yv�0����y֩NX��b*�`��<�x��	��>~�ɧB����$,*�r�܉����ú��ۗ8��O�ASL��s����Z}1k�F���t�ǿw�~KD��t���,nU�[-�c�Iԕ���G�|w7��I�+J���i#�&��5JH�5s��?4���nJQt��uqq����9�T��Nf��C��Ӳ?r/D>�V-�E�Ț%��d�N�3�C�� A��~��yFp�A��9��>f�,kEC.^xA����S�ݩ�&�0�i{�r\�x���ZX���) ��Y�!<�1=	A�s������^)f��u�Y2�K�p��Z�bl�������gB-�sr����!Q{Я^��ޫ?�P�L�'�[;�v��1>P�ѣl��л��Q�αv`���&���7؉���˱�{¶L=�r���zG�ϟ??�?W78��7�<�$����	�gY�\�qss�]ិW�Z��C�E앒��������F�ɣ/����,أ�G��t�Q� ��9i
V���\����C1��A^�k�$s�	QN���,n�Aq"ߖOEc� �k�1w'�@�
ӓ��d� �x�A<��mu=Z��ˈ�A�����:uvO��B��hZ?�:ԝ����m�Bg��;�}̄ǒ�Y{p�S�W6��:���N����4�ߢ>[���QbX�45�KXOZr;M���.U(.VT��K.�z�/t�0�`�@mO$����i�P]Z%��YM����6vQ�te�[e��)!�j+��O��gE��uII��]�/f�=]���9%!&�@9�Z�\͉>��*J!J�za����m(]�r���2B(yG?��c���6V^H��GBˤ(��yp����J���h�/��K�
Ry�!�5�Pv�tb>�R�O�YP��+�qm�,�!��Q�ns��/��I�:��K�n����;�O��~��7�̞m�B,A��"�}GPIU����8�@x^�o!�M�2���2r&&���('���Ŷ��R��'$t2��n����Q�8�i5��B9�)�i��@��(���+7���h�y\JHNOO�@�iT���9�`�\�\�/jӡo("��~�����k��2�����;�o��^?��8�A1�� �hv���w�vr��L��أr��_Rf)Tfv��"����]aP|������@ ��>���y�6��q�5E����[J��z0����o�z��H�/k�cG�P*�cN�p���ÏF�2{�0���5*����z���x��8!�O����xpᅻ&���3...J ϲ���>O�16xB8F�lO{��;$���o�#f�����ΨSk���.��Oz,R����������n�u�;�y����(3�-,@�bY�؏陙{ �:iF_�
��kQ&�E �X�ޛ�n�3�<�IR��"f�i�^���}�V��_��e�(�ZJ�	}Fʕ(�ѥ]�q���A�Z
���˸��QZ'Պ����7*�����l
. #�CAx���H���}�`W]�G�����O�
���ԝK����ҹ&��� �NO�'^�}��x4Y�n�B�syP����ҌVηF�=�q��ۛ�ڦ8�ߛ����l��_tL�F�L2��_n�����5?��`������4C��E-��y���l�껐u@�zt�r�O�b��F�i���Y� �����F�3-7{Z�����\	f���U��pv�_|,
�y�g�<�B~O���q����uH%x���\�Ȧ���*�ל�ڐ��Lby��U������k >%'o4"onz`�n5[;_�n^�0�L�uyyt�8���ߛ�����=IpR�j�K�(�ʮ������!25��R򍅩���h�>d����1i5R&�ht����7��7l�ZG�'�S���pjg,%h�8ǰ��6+	������ag����V�9;p�Y��Ly��,�����ݓ����,�Y�#�a`d<<ZS��	��P6�nL�e�e}L�>#�Û���p3G~G���Q�*6��+0�2(�D3�i����F�0�<k��<y�,�$� �X�呣�j�#�"���ޫ_j�T���K_�#p/6�ŻM �{n�݁{X#$����?�ﱏ^9:�Ⱥ+��r?��OD�ٟ������=��I��8dؖ�ާ?<7���>K]
�۝���z��7Ω�f�2�\{]��YK�c�� ��i���A¶y>L�ub�%�M�1VQnh��.Щ�DW������R��g&��-���>�z��5K$����qa���FIF�����j�_�<Jc��,�aN/���p���1��E��~O�a\3hO��D*��J�[��t6���>��L��V���p֚��Q���g��lR������X���]�m-����c�j�3���lw&x��nP����I���Ѫ�?�����_�u���k;�(%Y�����sbs�7r8Q���t ��P��B�զ���c<t���PҪ�ož�*,N����)����n��`�A�*���%)���3�)*KVr�E�h��W�\�=bz�h㽥��!HK��3���%��@)
1�u�wWz[E
X�L���8�&Ys#�1%uT���Z�˞��-G�5��|�5+�k�7�=#O�V�5«+_+�Szn����t�$WnG�<��Ep��V��D�;�T������7�3��U��J�C;ִ�/B��{@�����ܢ�vL���0�S���u�^�%}h@i�Tpy�S(
���$������
E�Ũ/��<- SR����f�qK)j/����/�T��Y���+*#�0��C��0e}ߴWs4u�(�s�&��B���Ɗ�єV;s��ot]l��(f�����z_m�-T�3]e���B�B�,�	7j�@��̀3**.����@��`d����� ����2.�Mǰ���>��6(�=�1Y�5!y:;�O>8�P~K������k��Q��@v����T��9���^%�z�-��4xY%��:� ��c<��ᑛ46��!c�;*�V���[��J���7>��ދ�ܿ��2w���h���u��7EGfS�IU�,���	u�t��?[8��<�b�zs���Z��p?~Y�jc#37/s�&ݘK�����ڴ"OZ<���C��q%�6x§s���5���{�
+��qI'�凞TVLD�'"b�nGF���g���\(�1X�Q�p�����,hS(���u�Л�P�*���[Z�hm}�CU@��-�^�Dڮ��ݓȋl��ǘreؤ"@���Y�r�������gi����.�(����}�G03����S��A���)t}�#��\��N}$����qd��5sz\[�����K	���Y�~�dU3b^G�� ���{?^]W�X�3���x����b@�;�k��J��&d@+F��$�#���&�C���� _�@�0u��8"P��ٷ�?���'�*�#`#��L&��	�ΪA6J�9� H�ğX��2���MYږvO$B�Y�'2�.C�;��Q:Uܣ���?pFm�d�h��ɗ��\���X�o�����p�!"��&Xwn�����&˹�Y%�0�`��)G9!X�h��C�[���_L�R�,�Гף��n}S'I��(�D�P�e�M[��]�e��:�5�����`R%D�cgVN�������Y{-pr��<�WC��sd?2�E���H�l�'���w�����c��:��^��fӺ1����y���p-9ߔd���D�z5�7�jQ&//V▩Ǧf��|U��9��Ƚ4`�ӗ�b����[o�S�������M����-s�[,WX����$��1\�!sz?��\�؅�Q�ϟw��"S���[
��u�9f��<g�8	��8r��r�ݖm�D����J�,b��%�+�v�8_Ё�}ű�ߓ���Н��Z�N��h�"*0:���ھ@�!�7�$;�:ǅ�H|c$�����r\����?��A���4N�E�&}nh�V7�>f���Z�̗L��� �C� 
�芧�FȪ�X�����c���'>���~��4~����M�X����#	p�c3õ���w���p%#Ƕ"7M�ьR������͐��x��j�]h}*��a4����l��P�}	�U/[����xS���12}��_�=��d��˧����1[�l.�5^+}�2�Q;�Ȅ��vl����:��׿�w�qϨ�z����ͪ�,�������;���X~K���T�R"l�_�OÓ�o�L���m_��9��b�v\�L�5�ҩ(� A�a���FU�{����\��O�N�=��p4&t�kK��N�%��Z!B��&VP�����tx��"�,��|���ʼ�m]�+��7�:�@�����C���u�oR��PvOZ����+� ��(��F���"U
� 8�)8/w� n��:lZ��	��VwJ�Mu��tY�mf�o���"�:I5]?�p-���H�E��g���eyK;S�w�x�SN�����^9���~���Go��A���b�����>zm����I0Y ���冿�H2%���M*�Ŏ���G����(�lOk���?`��"fu�8\�E��w?��t��c,�}w��A`�&1�&���\�~�G�r/����H�4!f t�4�H˒R��}@&q����ݎ�.�C�<f�ߕ])���(|1�	�1�$���8��2mq�s�}S��5F�J����V �U��m�����?��~oetmm������� �60��I�9'Z`\`����{κ"��{~���[��N�S��[ y����yI��U��!stK�����#)���Y�$��)�(.� ���%��*dF�\���2��'Ŧ��o�޿�0���!H-&��dڋ��Z]���`$J��_8��22�tiL�T|��_�_������ݥ��7�,n�o�Ϣ�� c�� ���ȸ�����'䖎�+Wq�A��}씰��?T�%^V�E���Vi8�w���ʠ${����]� �Tq-k��6{��1Kf(o���jOk�aaM��Hy͛m%���T�7�Ӻ�[pGa�����b�8G���}�o��XX�|�ú�+c�+�Bfy�>��N1��5O�,e<�%��hn��^7]�8z��x�2� [���x���T���oy.�K�|y4������Ϙ�.��]b-W�S� %]�do�g9V�{����N1�����Q2|e��3o������%� �7BXs	s~D�vy`��^���إ�Ҳ�e��ܘ3�{F�>���/��>=Yߜ%y����%=��Z �ƌ�=&����I�ܽ4����[����(��#'N3ÖK��ѣ���r��?�!���O��3�6̘2"�Cep��/�I	x�qvGv&�����K�犜��Z�� A�����^R析��t2�l��]�f�݇W���Y�{z���*�>YA�jΏ�~�V�o�lk5ӸO@�m�&���~k��g��/��f�SU�[aC=�~�o�'����k_��,�0UiҞv�o
�%e{�-b���W�k9E0��l7�9H���E�o��dR7�Z�@��9����w���(�&)�ft��P�����'���Fe�N�<i������1l��*D��MM��W�,�Nx33^d�4 ��[�6l[�l���ħdsqL��w~���f����'Wo��苆Z�N�&��,���$PH��^��ͻ�<���Ր���/#�R�0#����X�G9�ԫW�m�ug�4r0C�y[O��F4����4�9s�%�,����2Vh��I�t�����:�A���[_q�y����Gd:w?yG� >gA�d��v�Cw��! G�	<'U��:J�/Ѓ&)q�Ò�l|Y��mV6��T���~���yt��y������
	E�`└��Sb�FS-��T0g�M`���c�c��&���v�w.��,����b���̴�.�Ż<�_��S�`�?�C��k.A��Ϟ��
��B	��cIᘙ-��.��Zy	¹�f$����}�=��e��[����Ãe��÷UUU�����7���!242J��lq�hn�Ӻ���ly�`�9�?�a����y��筨�����"��b�����90�����J��[�7��������[1������y��@Rn�*��0�(|�z�/�i��LE�&�h_m�O�>:j�h6W�3=3}{Gǃ��Tn\�Sޤ����u����9����u�9|�|qd�|4�Z�!��z�[�=�y�kr�[���]ћT�?ۆ�����;��B���5��JI �d�
�=�7m�C&�!����＼�g>�揿�I$5Rb�/�y�����u���'o�!�n��q�|A�r��	o_�☲`n�880{[�'�o)+#��<��o�_�Ei	G;���n��}_i��q%x������ԃ��_v�x|y���G��K��Y�V$�f|�[��Q�u����v��ʔ�Ge����_�DCK���c��ż$���jlj�éc��H}���Я�׫����{����o=��yX��X(��{]\[]<F�w������SG����F*6�܋��[�~8CC/*QLW��m_aʥx�o�Bg!x����"?�����SR�H�oRgG������K����,�e��/*���;L����F����ˑ%���)K�<*���R�o�>��j��lo�V���Io��IYt�xp%f�ڴ '{#�%�"d��#JE-�5Jv܇\C�8y� ������D$�9y-��|J�����D�OG$E��n.�J���VzY��67mm5��6��SS;GG�&���]��.���1P� ����K%5�P�g���yg��QW'RS_o����R^Z�ty�1��Z�x�)�@��P������.��8A9 ����wB3�xg���A�|ځ �p��W���Ʊr��֮�Q�瞔�5�ߚ&�h9�!�E=P���vg�~_8]~�3�Ǽ23Q�y���n�!�ڧ1���y����$:&&�=C#�{���
�&�6�_G��>&l�M����{�p5=����v�j��z�[�g�&��Q�wr�(���aPe�����b�%܋!�T�KQO�0G�Ƥ�`���^v�Q��;G.C�c�y_��na��3<=g{�������TS=�444j�k"��PY�B�¬�p�����:��{�T9���p�o&-_?
�O��֖�I��k����o��˟��1?-H��1�ܷ�ߍ�2N����l��^��������%$V[DSK�d����|���"έI�9�?��Ӣ�iZ��W�E4�?+��'p3�y�[4�N�����»0J�j*����ɔ�O��{�z�I.T_Gcch�e�Z:7�v 5q�MGs#Ύ��DWـ�_eA5�z�7�f����Wv�%�8�(
�ׂ���t#�v4|}��(?(p���XA�-���>8]��ޜ�����>kY|M��m�<m��#m$���4�{�,^Y�̔��eE�sg��p�ͯ���{�����V#�sI7��7,�S'���Lہ΋��4��_e+/���H��_]�t�9�K�<g?+%|��\����Ua`1<ʯ
p0��9ğ�y�;��ʩO�*tǛ<88辣�8��;X�L4v��z��n��q�~v�K»i�C���$Zv�RS��P{rޏ]Yڿ[_D������'���[H�D��Q���G}���es����=z����676��2�fAߞ~�;�����!11ۼ��{�G������ȑ������:G�h㤠�!C�N6��W�^d|��֎���r{�//�܁555��ՁD��0�
���P��H
G��pi�pm��m�Rs�-��#QQ�bi��0�g������v���}�⠼�L��Y�-)�́��X�:N��ꣾe���*@�Q�'	�t)y:m�Zdü	m;�J)�b��U��g�jȪ��*��)W���-���?ƅ�� #Ejs�gz��j�����6�2��.���|�����G�B�p3�˭7�|��������//-$��`�"�u��|�)�n�,�]ˍ���G�PG�9�,��X;&���|݌�<ވ���2����ν��0L�R�2OW#& �ss���j`oَ��/��e��_:[��.��i%�z����������-��n����{\�ܭx��˸�G�ߪ�5�T���gf�����#c�Zh��z��S��keg׏v�U���]1%����>0W�ӗ�s���`5�j�*9�Ih)��^�[��|RdZG@���	��j��ׇ`���5&g~��^��[��u��X+��6�.D`�j�NlM4��6����H�O��P4�I0�+�a�.)TX�{22E���ھ�8��,sNJoI�,�W�|�w>� o}�X��i�Wo�+|i��H��k��5����!�<?�0��ͧr0 �d�e�06��	w:0@EM5�������|:p<��〮2�09������4 �[��B��P��V�ǝ���@��]�紿��|fKۓ%E���J�|oFH^35P ��=�iqC�H�G����ސ�VJ�;�l
v�8?(	��k^��<���s�,U;���8����S����HZ�?k'I<��檅��~OzoN���
��%I��3h�qO]:|ll�B2��H�����fpa#��w�y���"9)��&�4%+,��x�t�lxU�ҹi�8���	җ#��C��Ȣ���]n`z(��?�mo�	ò�£*�	�P�+!DVU̓�����'a�$�±����"�bn�L���y����_�.�u�e��ޓyΆԅC�_��M)$��h���u^�!.��!0qM���LF�0�� �TS�)�z�sű5�Y�D�{�����F�k'�i�X���_��xć 6��rź/2�#m��쮞�a�!!}ǡ��M��ݪ�-��TH��Z��;�P+؈_���䶋�8Q��#�8QQ��ُ΁?a	b5�_��e	H6.��?u�ם#�Sp:n��u
�yo�ݻ����*8��E)HP������)�-����+�q��"��ri�����M&�ZC}vQһ��e�?�����S�Y�w�O|������?BN�O�Q��¹�$]Jٵ�f�/˥�����9��+s֕g���G�u�C���J([ȦP���EHFF8;��l���PvI%�y�93�Ȏㆽ��-�������p���y������~�^�.0�7��N7�t�TE����8��?�Yp��ޝ����~�IL��'���wg�ݛ/�Th܃邟�"}<��N��Ê_�M�b�H��\��m$Dw&N�>���t!�7Bk��G�]s�zo����DQw��D;tO�+�5$T�A��/�ۏw;���
�{n�k�.���!<b�m�584� �c9�) '�l���
K�����<*�k{<㩙c&X7@[N�8%w�5n���vi0���:�����C���oF��I�S�3=��{�+j�=��OD����t90���qp+m�X~��lA"���:�y��ݙ�!�sF��_*u{8��gu�*]W� aY�7|V�u�"�S7��CL���^�Q�O�>���,�~�'ާ��dgm�3�+�fVV�}.���O�);YӉ'ȿɀ3�;�wr�md	�̷cy$6���(��~oj�&���Ϙ8���|��.)kOK�m]�$KH2�Һ�nv.���i#���%��fb����srU$�i�R3o��~!��7���P�K�y�d��U�:zs���~���/R��v���:�X�A2�B�ٹ 2]">6��ٌ&bd|+W%�Jbbbq�˳ Kl@�T�{
�%ꅆ�Ʒ�P���_��`�*b�[?���(EQ1qm��[���R*�a-�~���<[&3qa�q�9H��m������s���;V �N��fu=��=o��3��%����1�ئh��LȊ�VB�b��I5�:�${(�*�{�ݫ��N$θ�q��+S�@���n�㌑Q�������j�/Z@��|.1,���.����-�y�F�3�H�����������mCE����dM�yܴ��7���Z�]�D<?��M��Z����e�JN�u��>6��(�ǻ��6ҊJ���Uq�g��oS���bb$��Q�]Vv��^OZJ*�7KB^bb8��}�e�3����ܣˑg^���SԤ39{��ki�o�_9B�B��8^>�j3淍2n�{����N��������m�Ý��t ���>�QB����_׆���SWpo^x�d�5fl� �"����#�̞_zd���&�;�Ւ�j@^ �9���ύ׀Y���"����򮠠�$������YV���W+�R����_��TUk>{�K�3z�U0�`�ڧ��6�f~�a�˾A$�W)��\T=������U���'�jc'L���]7V�A���}� ��%ր����`!V�h[���_�dq���Fɜ���z�r'��B�R�4�>�
��W3�1p#?�\W���rX��8h���P&�?��^K�����~�K?�7h|����D�nd�8��?e�cOR0#��2�����k�B�+�G{�uc���CJJI��	������������Z��>x�e�Qڕ��g�SOa��X6J���;����K,�9<���ҍ�߈b�x�������'(��ƷŁD���������T�mD��>){[�L����������w��{��&�F�/��R�;ż�iu�k�&����߉%;�w�siǮ�^�}Y��޹�}K+\��T2J ��IsU0ݴ9}v���e�fO����T��3+��Q=��X�0�2��5.� 6��Y�ҸM��q+� 7�*o�T���<Q�+�;e����`��?u��?L0�v�ػI��b�zy�dqu��C�%�.��>�/	=~'�T�6x[ǐKB�KU��Sv����[�q)�nzo����K|��m�8����R�`�̔��:` 1��I� V>�P�ȥ���:�| �d���Q1Z�2�u�2T�,99�,�-��l`��t*�"���t��~r���V��D���?Y2�:�^3��q��aQ]�I�Uy�?�F�{q���wl-�_s>:��V�_u����ڗ�0-�gϤ�u\&�(q87���R�H�rv~dd�?D�WJ�D�I~��΂�O� h�>�T�$uU�6�x�	/���� G-U��$�R~��z����<e����򹌆�
Z�'�n7�b5޿x�ٰS�@@��&m(AH�r [�{�� �3�9E!����B�E�_�1�wޑ���Β+r�8��`}tR7��͐v���`�o��Ԁ��t���G����tRi�8�#�(����t��ژ�J��')��.���:�
qzwy!q9z?o��C���O��'������D9�������>�����r�����T��Df�G:���s鹒ᱺ̱�Ci.���=H����xT^4�����,s..���-�k[%7�Vs��џ��L��ߕ�� �������t����6��HN��T��$�V�v�]o�ǡEX�#�R�]/0��GKMET�CV8�^�)|���|X��^�����xA��~G֣D�&� �.p��t	_�f؂��WVA�^���Є+�K�ܖU�i;^ի�1QSS_��P���#^��
e�_�jh�W0������l�z�`�h,+N'QV���V���';�n0����l
��~�f��V�#+r��3i�g��m�_�?L(��T�`�]t�j|/K�����z����r�Y���eF��f�l�gJ(����6�;;'gs��[�W;	4.�[7D�6�|���X����8zI�AȐ^���qo�N#���ys�ٞ�MT�퓿�x�C�xi@��ôz޽����ф��Q�X�Yէ�<J����F�?�����*�����j��W����Qɏj@O�p�
�	�\}1f��Q8�Q�r��ǩ���דy�)o�C�-�3�u��A�U��ؑRWO�e����č_�>��M�Pz�-w���ޕR��N�Z����Q�^�x�Xkֵ�|�]ҭ���,;/(y�+��������,������(�N��6�6�_��ɏY�eNI{���ֹ�+�(��y"l*l�"W5���$�fy�s��[��m�}��xA�����x¼��唶l��k�׹?;���+T����N>5��%���)O�l��g;F��5�x�u����[݋F�ͺ�	�T
�D˲m��uu_�wn&�QG�˅Gu�\�q���b���M���j'1��܁�YK��ҩ��'a�^��^G3.����������r��������A���2���eWq3F�/j@�V�����!�Q�^�����9	XA���QO?�-����X��bZ���U-��r�?.��{�=]f�)���sn^��k۫EGr&���M��<6l�4��kW)3+���ڇ��4�r�6��b��}� �;lY�yݻ���<�^T��^TkVҝG9:!bVL�?��V�-��K��v�`�ԍ��ŉ7)��}6i�J�@>�]5��c4�ː5���tw%fx�JD ��0BXb�N����V�I5tka���'ğ��\C�RG��ϡ�G��0�����/�[b��K����	'��\�R�����������D�,q��l�7o<C�3:+�X����2=�`�-��Gu��|��Pvx��t��(���x�]������⧟¾�4�J��|2��Y�o���T�#��/cK�?qy�s{�mA~�i���q�i{�;I�t�ƀGAn���>nE�����仩�o?��xM14�R�*ȽI�K��|V?U:.��O��8��3?k�}9�X�r�ܡ��K�t�?[�h�U>�~�bp�i�Q܇z�rq���n_��:B�G�M� ��=�B�&�b��f��.����QCp�G�Rr����@UC`�䶖�k)�KwJ3&sa�X3�]_z�y/$��7m�R��2�jd�)h���Ae��(~q̐=�w���|����پ� 0���a!��I���O�,t�j��SQsHTO�����E����|#g��1|=��������?UԱF�6,�x��|V��5�oWď�+�N{C�O ��"""��3��G�vI,\zO<�\��~N����+6����_����N�R*Gm&ښTJxtp�0�����������ALej��4��\��N�Vo���鄚�r\��fC�--�~�ao!m�u�m���JK[��� ���q���iJ�,���?�3<`rtr@⣗�C~[ZZJ ��W�V����&�u卦8���!���Z��@~L�[�]�;b�s4���n��ė0b��������NU�_r�8�+1����Q��\�5��X�kUp2���"�m�{b>�V"������p4k�?t��B�P��+դ�Dt�4n��`���(�Л��Q*Ȧ��ײ�A	\��p�@�������W�<���w�4���ͽ֌Pb�G��������S@$����k�垺K�u��[}Ɲ�i�&�u�3?������'����(��
�z~BOAZK�[)�"J��[xL��I���s�,i ������������T�����<U�ҋ��Ї��V����dϐ*r��&4;;�junD����Ld8\�jPB���v�A�+���u"|hA��gE������7Aao1�>Z��!�+>����L�f/)K�=v�!�AJ��O���,�W�p�T����`SV�b�R
�_>l�f�{��'?5M� i�����_�Ik��+�B9:����3�1���<�$8\�������=X�ͯ�����P�-�m�W-�D�6��@�g�<���𖯺c����?G�,��?%���V�"{Ž6̺#rQ��yq����(S�Χpé_bO4g����*OlC"8c��Q���!�j��;��1E��*��\h���[5B����L
�{���e��а�I���˾�*j���(:O�7�,��I*�{*�R �d����͏r��R�nk�e����4����	��QX�=�E{U��7��j��.��'����@/ؙ�K�Լk�"E��Z��
�;�G"w0�}1�0h�:V:!�a���c�_�&����cep�8��՛���2kh�[]___�T�a�Q�N��bl� ���h���i�q�о�m�:1��d��k�����[/2ֿ�`\���+�A��A(�M~�
D��j������
.��O��e�����Ԋ.8w��睇�!Q`�g/���ppe�G6����F[��6������m�6�Q��Pg�:��o==T$s��ML��.g�½!�7�:�	�M+x訾'oUxk�N���I�".�/O'm	ǣ��m��=�
_�]Ѫ�{o1�+H�~�V�Yո�[��z�:8��
���:�-�}[���+M�s�ᣛ��i*G�˓�;��Z�%w�����Y�-3'��~8 ���J��0\��ڞ�E�&� �KNu�8b"�����ٻj����eK�"��yߑ��;4�{�w�?�v�����684�F�q�9�e_v(<&��>�B����IY̛!p5<,��,˳i�=�#��o|{4 ��ZAu�jbw��N��$�����^�����G�T��h{�1	���I�UXt���G3:�Zj�[[���ђQ�cM^_�QTZ���TT�����j룇&-ˎ����{��U�ؕ-;����m�d�7��W��F�.��UA��.��͑�� ��D\ϾƠ�[:5=���  �Α��`e��w� ��C�o?zI�P��M�r�[��D��˦�۳�$��8w���Y���n@_h�rXIԓ�έ;ƃ��w26c�Ėdܤ������Q�+��Ӫ���_�D���-o��>� ���t������&.��``?��-�h�Zb��s-CԀ$�X:\��P'�\����#�|����D��)��zz�SU���j� ��`��t��i_���LF����8�G����߯q�s�;r�^yNP�ӸR� ���q��z�����mm<c��,_�Q����c�F{����y_>(�s�<����l̎'j����TҸ���&#>�a�I���C��^��~����r:S����[ uL��~A`F��		�z��7���U�Ŧg��7K��PP�����f��H�q�j��I@m
{�1���ۍ1���X���&�q�϶�$1��j���L�
������J���Ι��by0B[n��&��>�,�E"�>�4ݙ�6GCwg�tXϲ
�)=xÙ �X�e�Vt�����1�Kךm@��:�xVv.ޛ�#����������D�v�W[6� ?pj�%�v6.��žVdzS^s{�8�𫨷)�ŀ��);����Vt{ښe��e�W��T_1�,�D�Iɳ]ץ<�}�z�����1;��¦�T^u�C���w����J(|_n;���B����F�n�j����đC<�>)���G�u�W&#�2qlT��:
�ꁷ��\ݦu �kB��ҋ���q���mQf'��ٔ�'�5`�/�3��Հ�1����kx>'�����5���;0v¹]|��<�/&U��}�۶��:���]�������0�A�������y]�_���,G�=����D���6�����d�A�55u��B���Ə�+����m>|�pitq��cؚ]���1���GH�y���ε5���<�=E-�;�|���\��yb&��N�����tS��:�ӡa^\ǫy���[�9@�#}7�¶')��:���1��&�\�}z(*&����Q��\ɾ���cd�s&I���\ӯ� ��w�����&1��^y��;Ys��v=ֈ�ҹJH���?������F}��]Ϟ=�c�%a�I��FvvN%x`����ҭ��1p>wSVO��{Uu=�u!�Սj���%������iP���_��bjZls�B��(.G0�.�zU-Yx����{"r����]�Vlv0VN��y4����d^D5V�8�&���hz��tѵ"�c�_��c��
<���\8�4�>��3b������%OU���kmi����.�?�r�d�&���@6V]gy���v��g��F�~��@����l���V"�)4��gt�qoHws�D�i�L{�TM���#:�ڼo�ρ��z	lJ�[_熽h��7SݩҗSE�Ӥ�wf����[��x~���v��9�P^�`}S�jZ�hD�i���JF�E�C^����٤�����h^����*K�q[e^+v��߷E�!V֋���߸?NW��f�G�W�7q��gg\�dK���9��W���v�u�^׆�~�2�^c���OW�M3�lM�m�(�
�P�V64��E|r8􊮘��!��E�΍_K)L���b	�Xn���f����?#U5�Q11�"iR&%r%��>�,�m�nF�ش=sI��y{P�������CR���{ͨߒ�1/���P������8�j�G�k.�� �2;�U8���;nw��z������'��1�aP�P���#����)�kn���$>��(�rk%�r�鋆(�>}��5וL�3wV���;{�/c`�֥����� A-�{�ޛ~���ٕ��	��8���������ɔ� �[�qq�������^�;�m@�K⧭xK	j7`��q�\w�r�q��)Ks�-�Z���a1ٝӜޤf;7i������\�M��ĩ̴�L����q9o���6�m�<i}��_pSS���b���Y��~�'e7=w���^)y�ߜT;��h���
R&�=�/�d���D���߁�%�g#����F�T�������V��k�m2D�%�fQ�_%���m:s]ù��K��)����zzzU[�?GG��#Nwu"�,G�{6�O�{�� T�j9|������y>�ϔO�&�!�o榇�7��E�(5 ��Yvw��@���I��;_58vb�]F^�l\F��2��Y���@��d[�{�'3��i�un���M׎�r(�֬�w2N�^U�=�n0ڦ&3-������1KGҟݹ�.��N��1���/�2c����=b�o�S.�|pa _U�����J���՛͵}��]S�g�|7ȏ��7���1�T�������m��ӯ_n^�����x����5����ޣ<~��7��칺ۿ�>��m��u�����ډ��7�1�d掫g<2`�KI.�U�y�z�T֫����`�?������;���ƪPBS���	.X���5��$��5G�fƭ,����@���0�i��h��T��ȕ�b�j���p{�2ngLy�1G q��	�^�P}�|f���J�:�j��qX������*R�Y�K	��r�[R�<>���"M��a�O\��Q/'/�R�����Kq'e�4>s ]D���-���3119�X�W��37��l�rX\⋀����ܞ�KߩJ�蕭4s&UHz�]AR"�/l�`ط������çR=.c�ymmm����i]c��M��珛�9��wq�=�p�%%�B��8�<��2O�� h��]�`.�<P^��,�ţ�W���H�ұϴ�l=�]�a{��S���sx!���IZ�7(����������#/CKf���K��-�k�~(��8{A�H|]Q>�:�RTCV���Xq�,O]511������̲�������.�Wn�	Q��v��G���h$�\F�h�=ijj�z`�|W]]=U�fz�>6���W�!\ⓣ�OAN���bf||jT79���-�C�d ������]7��Iu+����:�vX�"��>�B�����1�)�h�����|�ΝS@l��Ċ�G���i@�������mQ��Tju#��4x���P4�4�:�K=��0mV���u����M�z��?Hdk���l-�,��eKe1K��ҁ߫l�Z���� UD<�&lߍ`L��,u -Ҍq�Q����	�TaS��ȫJ��=�?�_�,��f�����a�dWkv�ڎ�A���ч t'n�9ȜR^i>z��(�Y!uԀ�n�$�`mr�J��gl����I�X��f �}��H¤|�p�����^\��g�K���!��k�/�\��L���Xb�_2 ���]ȨϽ�̴9���@}�w��M.133�;!6XX��C��Dk5L�!�ԯ3H.G.��l[2�/�2p5��D��U�VەURV.�,B���1����'O�e_����L���Z7ZG8��p[饐�����Z���t�lF���O/W��0S��v|!.S�1���E�!L�d��Ɏ�<Wh��kk�����w`;'���K�Ye`�?��D&f�e�	.��Q��@w�/1���,OE�W�JW�!�-g'O�<U?����;]f�K"��CH�uׅ��h}�=i��l����V��.�x�[8��۽��e�.�D������%��� ����}Z�-���2�4�B����|��j�`�Օߕ��g���>|h83�Q�2����ٰ��v���꧹��jr=��J0��R�l�������/--=���6y�|�JfVV����r����W�x��Ek!�����?EN>�ʞY�fe������}�V��d��7]�tؤ�G�N�ɠ�N�?���2�nI��ޣ>S�dd|=�pu�z�����5���}���O�uu�jjj:���,��vU��E�$����'������#�$�������x{jû|��o���f+�p��:���,5�����s�MA,"��w��_�}w�����d	�S��}�w.�=���l�H�Z&"�����d�~���}������%�:y�B���~0�y��(tL\�qZ^Y�x8"�E�!�~��,�(Y�o�cn:	u՗��Td�nmI,���57�����9{x���Q������EB����˟�����(8[�[��A�豱��|�)�� V�����AEN���,?���O ����=�8�&�4�ɞ~�:8���qΊ��cà��i��[���,xg.��x)n�����%�}ڵֵ<u�r�;�WJ��`��l�Z*��"�$�����3S�΂�#�F����̬ �־~\�JKf�k�w�����p��p=?Ԅ�#���O�Q�M)��h���#��"�=׈~�N�|������V��d�lg����*���ٿ�f�_�;�Lm���v���A<	�����uz(�M�W��$�T��o�o����#�55q{p�Ş�k���ZG�@%����!��,w� �
��� ��a]����H����)���T^{,2���������m6.����l���#�SZ�M��0?;������۽8�=i	��"ps;���g;:R�����!԰( �W緁�1��oTH����Q?�|V[�x�ؾ�C�;���CEM�GA���3G�>���CD���ڹ��ǚ��1�"�����U$���we0�+!�ّ��HnTG����O�\�u����]��;�����Ilf/���@T���_rAt*�d�X7u�8�P�1{�r"���҃|�+k��l��\���EMd1��C���������ײ�rt<:�TwZ��B΄�Uq�IڠL窈��(�t)�:/Z�j�pJ9��j��ׂ�¬������K��b5��VxE'#r����84�5���]�L��Q���4Il�p9󅊓Y��T9��w�����t�)�#m��;�;<&�L%|xH�����Cv&)I�mv�gjXa7]��1=��#�l�±o7� �sX��&M���C�ޑx��c��WY��5�ޏR�7m%id��
�!�_kVA�4׉��,��]�u�R�@{�I���x����8,lI~9z��^]qp�$�ͣ���78o�����d����g��Pj�
�K�D�}pg� ��X�"�lr�"_Ѣm�韴T#d��KA/fI�.�|6&Ue�r��%.�T�Ti s�C!���w��t�>�x� ^f��
XK����.'��ܢN��Ng����%��r��n��G����O�U�u��Ύ���e��|�JUg���gz�:����l@����ظx4�:�u��%yB�!.�R��J��T���
�%p�w���e  �i��(Պ�CS$������U�Wu(jn�oܨB�5����Г#�	+�k�������P��wo�(��)��d�jW�x�?�[�6���=cZ
!���F8}��H�=���TO�'$2�z���*����?�VA��@h�C���c@�{oRܝL�۲[�<L��[�譊��E �VL��Up͡� ���d�RS��*#�>@�o"8�t_��1���_�wxr{�@���GY-E�N`j9����N�|��_����Bk���A$t|�j���v���W"�2N��sﭏ��{l��|Drܛ7oznL6�~��:p݌�����A���^J=�;w����+*&�z��f܇���i�����QI�r=(�3�#}Mxؕ���$eh��(����fQ�,��%�ث.�Ш�,��=~�AW���B!�{Y��)k6_<Α��[�ML<�oʿ��ɓ<����	c��>k��m"�KLL�M9H�1��r��P��/X��?2��mq��_�/T0���������WS��i�Ke)_T�X�� o{�.�"�>�Uz�T�U��x��i������#|�N�<���w��{w���8���e�b��pA�.3[���h�����j�k�F14F	 �4;+�<�ya�cV|�%�$N�!Hq�լ>r1��#G�J@ȵﮡ�w��l"B%��^��W*��P�z1Dqt�>F�[����/pT�_���n]B^ N��1!�T	�1R5bbD~-�ލ��j���Ji�Ԟ���C��KX7��"��<�[$���XZ����z�����ݽ�x���vu}*����h,�u����+b���aϸH�i��A;�|R@AO����z��|��O.�ǀ���
��N���N*8�/�����ܔ��}�/�؏�y�n�E.[v�M:,�&���`k�m�k��K���T8�'W����62q�Բ���tB��]���^��>��I�(HT{i�aib����Kc'�Ͻ����j��c��i�<��A���ҷ���ڌ�_�``�_+̻�d.^�1n;� �m��q����TC�,�k&,"��u�������ǒ�`j�5L���[�$ p�^�,Q��
�b�{�F7:ÄVG�_�ɴe0����x���d.��]W�f�#�2��;���,�$.'����@g;�q-��cء��2yڕ���#KgR7�����&�)�%u/���(S�{Lv����l.��y"��T�o���8�x���MpPA29Q��M��>K�����'��u���O	�K@��
}�;~V.�*@>���G����u�'bY��zC��.϶"�(��+M���B{"w^��V�A���KR��)\�ŉ�w�s>��+�.�n|�nBE��'5ϸ�D���8d��a(��IC�|5@��:G���C��.�O䟬�	=1b�Z�0��' �B��s�wԧ�{�����"#����%���qe�q d_4���g��m ���׏��޲R	�)C1�1_��f���r:;;z����U��%>?��zL�bD��h���bMLLd[���3��;�P{���8��<}�����R� \��`���c2�:��?�4�"ʽ�Bt������u_�3���w��ܛ����xo�*��m�WI`�����ﾸ����W?��X�Y(Y���e@/��yo��S�����vޤ�� ���8�q2��-��=����t篡;ھ.G2��u�o�'�>qr.����k�	ۚ�e�ݵK�s�6yް����%�� }E��ؚ�se)Q��~Y��<ʟ/��/o����5^C?�����E��~sc\�=�dt���5��}-p[������(���]�d��A��<,���W}��xh��q�4��]�aF�y�<�|�"�́!�c?����1	�ac���MGfq$�7
D���-�,�W���jk_!Z�a��p��}�˓=;d��W3N�����9����v{Y!3ߢȸp(�:<��\�|�ߺ�"i�&?�zo����z�i3�WXޤ��U�:��-gj27	�s��
5N���ͺuX���ҲM��r-��
BRv��Vʉl,�6��&�����>�У+��̼?ނ&�`#>�؟���||���x�ΐK�U�6��ߨ���T��U�y�m����郘E�&b��3�����qi�e�������_�s�c�>5���>�x�G�i���|AҒ*ш�}�M���ܣ��YA�*�9z�h$��
6�QO��P�s�=xF;�)�ؽ��D�5�{��������P�ˠk��P�;RO��b��=��[���Y|@*+��?�AG��ׇ� '26b��S�znF������A��:MC�ȗ��2'���9���J�繋��1�.aKo�^;Gڋ���șF71ӑ&���'$���W���|�����h�7�coM(�p�[��H��W	=���i�g}�C��D�O�������v�'e���s�jTLw�ܴ�<+�G�E�1,�A^�=O�߂�^"�MV�?�7�&��.Ad \���/�$��Q�eD�s��&s�#8;�0!�V嗫b�e��p��Sz�ެ���)��L�ʋ���wz�=�T������U1�6w{y�]Z���d�n��D��g�r0{����?k�q��ۄW��Y~ N����О�Xu�n��i��	oIy��r�.����/�^<=~��+A�J�_�	�����{�G0�'����۴j\��3��6O�$����& ��Z�7p�,����1��2���9�Jq�7*[���� uѷ	s�R�|D����M�1O~t� ��<� M/�w�+�&=�!�ܽ�|5�7��J�a~�������\���<�p����m�,������fy�ٗ��$k�h���D�[����4��������$C<�UO����m@�u���u}t�<�e�����"�Z	7~xm/0S��c�@��&܍�B�<���%�.�p�?����"�A7�9��m�:ٹl����C���te�4hkA�����2�jw�����)�f�����ku����&�l0� d{�����se�wy(�����m6�v.��.��l3��v<FkN4==�>���� ��9셍���b��h�n��/���q--�|�r�D�â��z�D�q5�0c�d��/�<�K�*���ᴩ4�8�"���@XcA�<p�3C���0��3iqx�IsE�g�A�#�ר���(�i���S��������g���I�1��m��A�_�`�klJ�㦌K�l��70�Y�h1�X2���^ƬX]��=�5d$3j�0c���hӿ��ၽ=�"�C��C�h�h�	Ԭ:���嘣KKKe���g�O#l�.�����SR0 0��g�Я�l��LRg��(yˮcH����,F��i���Z�q��;d�b����<����n���s�ܡ&PP�8�F=��k��o��p2{��]�E]��	�����G7 (1��{i6���_:X�'��䙥�u/�#x`��z�߇o��W������~�;�Rjz|�ֲJR���((-YS�e� b�]�*��/�Ik�n��j8����^���14:Q룜�� ���Ǫ�N���������b,]�1,��#����yӊ5�}_���U���3�K��?S�j	���Ls:"�y�0 nk�E��܂��X�T� o���P�7��p�a�T�SN��N��=�>�Vf4|4a�����L���&��J�86��%�8�)�I���-���y���<��֤�i�0�Y��@��^����u���2��8�<��x��)�rD���e��.�`t���\�$ڏ��T[8�^������7�V3첽������ruNZ:����CM���[�[���cEi&h�"�wê����R�@��uh1�a���7��\p��묢�;&<����G[�W���9ý�u�����d|!]��i꺹r��YGiN��^.�������[,���|<�ɵ���e)��V>��u�v��_��W�GQ�3E���r�
���d9����m�N��n�z����z48v!�}Te�pB���D��=�z2{'P�*R0����B�.JݺAUa�3?�V��
������DP�[��^g��X:�ΰĢ�Mzu�/��ͳ�G߅Xb�V-�UC8Ƥ�#eoOSqkR�1˻��X�?������5���<4�l���v�4��b�'� tvnn��RȜ*�7;܇Q]��~� �b����䛰5;�
�����x~��l$t�T���$��5��坖uI���@'Q:����l�ʴv�_�ت�.0�f�j�@^�o�m�.$<}��%��y�Ȩi�T&!���-�J@սT�D���I
�FL�T7+��'�-ɽoU��F�樨G$ O))�=��~/$Z1hM`������D��P�����2����4���;p�[��{�g����A>1�=i��ۉ7�iFL9�C!���̞Yj�P�5e��L�F�������-���Pn�Nx�GL0���}��5L+mn����x|íb��;K�D2�Ġ�p������F_�Ah��'w_�����Z�T;�������,�8X�,�>p�iY���7n�i�/7??@�t�a*!�P!5�p�׼Bs��?��s�jNf�ϕ�� ��Ƈ�9��X�� L0�J�6�F�����rmu׉g~��"�7R(���nhDۑ/g���dH�@�)#H�;���k݉��_U(����n��'M]��a����]^��'_��R�M��#������]t}��aC�hzz c?
�_�wXH^�.�ዂ_�9��D.l�J@>�/�}ت�V�4L�U�=j3$��&T��,t�ѹ�o���[9֝.��/w�U;�v��s�b=8[�♜7��Q?V	��W�U�Y�ZP�x|��������������?��q�����>��Nc9q����sݜj����IU󳊆�D��	�]eQ6�,x��6fLc�j4�/i |>ln���D�aؒ�l�����J��1a�Tˀ�����Y�*Θ�ʾ��m�^Jhh���H�詈�d�j��O�����R��K��g"h���s;�i0}��u���>z�W�*�H�Ɲ'����h�s�o?����^��@*�%�E�{_��mddem}�&�o���4���YW_*�<iP�v�+���o�"Eg�)E���M����KY�=��?��R&�4"}d{�����7��V��c���(��K�������l2���d'g\* ���)mU�Z ~�����VA����;�Ʌ;3#��
�s��&�����\t� �q��Ș-PX�|���ѝ"��ՙ5�ض��ԟ��%N�뜞|� �u�x���D�d�����Go������	�������{�����5*bz8�eb���R"�0ziQu�����0�Q��b��H�͓�������.��k]u��ǝu�KW���]f~����Έa��tI�fq�'��/+����&����q�44�׳z' ��mUf����0W���!�z[
�H̙��.w��d\���#�>���JJO��xlO���Z\��cߞL𤐽{����W����f���(^ߚ�<��vH-/+���$��n���[�la{�o��{���%r�OY�?�v|�F�?I{�B�;~ ���[ѭ�q��&�4�o��YjF���g��S�r���Z�$��P�2�Շ8Xji��1IvĿ��67Q�t��ͻ6���͓D����V��ǭ;��E4�S.ww�i��?,�Xv�V�*0em���uu�'��}��*� E��!Y�N$X�#+:�=�F0D�K@r�I�Qr�#���pw|K@�Ge�����x�����(!��E�M�3D*#YWF��q�k${��ɾ�.�ȺHH��^��6���5��V����xxؗ�=�s��u��uYm��A�|jt����D~��ƛ����ƃ�\~�'�|JP5��6s�����7��Z�/ �d��]8���9!H����i�'����)ke���	N��y�_r�&�6�֭�mD��zд���=P���\�ᾱ���ǈ�P�ڥ'a��ͭ�`D�_�4#7g<�i��?`-��}a5��>�YO@7����<\���3lMm��`��S���*��IZ�6��8����W��ԉ�l?�	�^g�Ҫ�V�����H�ݙ��sÅZ𑉷1�S�
6���}<����O���R9����FJX;��L����bV��ٚ:�/xM�������M�|t"{���gb&S���te�Ѯ�P��������	B��,a%���<��)Hp@���~<���u�����NR$g���n :��4���bT햹�2�+5�'��~/�d��~��E��
ka�Z">�[����3z)��:ŪkgG�Q�-<�J^]ݽ0*��,��w�����q?b������}ݣ�[�nǾ݆i
j�J��+�%7ا�����Qv0�~~��+Z$j�p,����H�}�zs ���p��f�K����޽E���cF�{"���?�>�\�?C��5�X'�%Fl*���7>|�A�*��ھ�G���������O����Y�:N�i��;o�4�F;@IJ��򒪊	��s�
��	��z����y������״�e��h���f��FFc�N_���fV�~l�me'<���Q�qs�JE�༎x�[ )�1,����ZgbW;U^�1V�Q��H��8�S%�i*|�'�����eC�G�P�p�5�?��Tz��-:6L�UT�;	S�;�۱��)���=�D@�ږ�`���n�-����ȁ-8�:�܋u���~U{s�k�����NA����V'\�U�w�uL%�yLF+ϋg!"q���7�Ŀ�0E��U��uߴ�}��염���vOZ\@o���~�ư6����r9�HzT���k��9����D�I�N�34��-���8��N��NDT���HT9@��&�+ۋ�̧|���Z�H`ܓ�#���-���x
-�b��D�I`�6��{�B	�K����I�3�����^`)-8t����6(�E%�29y�OD������U5�~*RI�RG�	�w�6�$=�&2x�pKp�ޙ�24r8eLz��5�U3Myp�x���x�g�������F�B`�Sr��Iu=�fE�ӗ�I�'�����>���� ��9IK�g��y��6̜b<ot14xϘ��C�[ �Jbr[j`���S9�ן8\�aY�Nֿ�;j���[ ��=�\,�>kx'QtZ������|�;�u�
�R;~�Xo�[����K�"p��b8KMH<���)�K�����|����%���+�Gx.�&�����������zߑ�D�n��`0;���{э�?���F�TLY�_׈�v���>`y�W�������N��:3��/D�7U�_�n[b��zj�RA�g�F�����~���]�)�ϵ��*	l�da~an��7�hTy��^�g6����2xn˸
'im�����a'i���3g�e���`��͖U����$�((ɠ�r��S���U	.ٯA�b�6g����/8�9|���ǫ��n�%�7��9s;�u����V5cj�~��$��R�3B�V8���{�éhu������c�掤O�=��~��o]&�p�'�:H�{�ǡCM�IF?�0u�>]�����47�mG[ݎ��^k�>�UJ�������+ˋ�mǢ��z��q����oC�����v���jfEܽ�+�=���|�у��^��_#z��ܚl�Q��Ͽ���x
9^��� �^����V��gNI	w��ಌ�3�NDssW������2(k��� �i}���_�sC0r���y��� �d��~�5*���1i~�+u0������ s�ݴ=1��u]�z_�OD�s�Q0�y��n����ln��e܊�t���zI�#�~�$�k�g>�� t��ڂ�P9�J~�́Ć�h�2��lFcS������&��c[��.�G�Y��z⹀�Ŏ;�k ���o.�� �l�-�(��d�Q�y�ȕ���7Y�1;�:+&���k�"�V���z{�T�hJ��,{Ȓ�F��1i�,I��Z�~����0tmn��H�T�QϠ�2������e^�m}��V�B3�#�r�1$i�ۡ�=C,!Α���ځ��p���7���ƛT�S0�XS�����*} "���f1j����=@zA��p�P�������:�ܼ6����}VW�ɲR�S�u8r�7/f
���M�	Y�Z�B�ùT۸�C�~�%�Uܙ
���ݾV�v*�l\��G���?U_n����pV�]�LW��y�p�6�y�3��TGֳغ�������}V'�b�=������ ے^��vV���q���F�9\=]��Ǜ���:��*�m!턶u�m`\x�^�s�J��k
}Ѵ�Vɹ����>Ҹe>fW�t/��6`��^U77+�z�DMMmKH� Q���)�n��2m/_;�?��Ư�hٴ�zr���f���嚪��6fe�c	������c9}�O���d������	��P�1�B�U��Л9�Vg�����*  ��K�k�����BTTT_p�'�+�R���+~���+�>�Z���~�*..�/۱��m��-,�L�"��z
�D�5ɪ�h5 _q�+//?�����N�ş��̍gc,�认��CwQrq�q��Q���)�t[��)nf����f2���3^��m��UNp*|�^?��qb�CÛ5g��.���i�c��"~ Bt\��B�I�Ґ��V�_��u�֚j���Ό6�)�W��Ln%j�/%DEC�v��n�͐F���$�.����}sf\b����
3�9�[R���5A����$���GMVI�N���-+�B
�S8y'NNI��z�
<�p�����-���?�N��S9�v��uf�D�;lλ�o5�7�R=~5��
?gH-�8BM�qs�Ip�-����v��Ru�Q���cdB�A os��5]��ocI^7�Zgٞ��V�=��S��:����˛�Ξ�}��+����2$�#�gK�m�~��U��2�J��GU�0��:�����J]����M�2�<��؄�G)���Š��3ζ���BWשX���l�m�=�2=$�K��������@?�V?�m��~Rv�{'B'm�9؜i�!sn�@0U8p�dacc#�B�É*�����l̧	�}����������ߗX6�
�^�����1�R����#�W�9���`��Q��>�=#*��X�c>�x�����b+��E�+�<�:�<0���@;�ug�*��싞�����l�:\[��h�8�d��v�K7t�<\�A>��i6d��q��$]Ӻ�s������J*ԋ���ܹ��d�=]���.�jv,��%]sY����C������q��B�l	���sQ�K�9ʹ%.<u��������Qr��4)B�v��=���n+{��&��2��7m�L�m�3b�ʶń"�E������Sљ��AZZ����z�ӊ����DYTLlع��׌��羅������!c�Y��������jDsHp�:a|����8�������RX��y��́�'Y��Y#'�"?��͔��4�*��x��6݆�I���RYYy���8�tB�����M��v5rI�4��yi��7�_f,y_�/<}Qy�
շ��j�`�׈�/�{��s��9R&{�g]��t)�W&�ʎ
U<@tF�Z�o�4e�!�����nK ��e*_���8�(#���*N<_5S�����g��|����X����G���r��*!^n~O��/�iw���T�'���2�e�pu�fU8��7c�Z��S���=�O��!	��E�S~e �j�͎�OZ�w*���vǣY�=�Y��	Wם��f����IZ�1K�A۪���;�n���Dz���e��ñ[��c����Ӻ� ֺ���S���ӷs�(�3���*߾�da�]�m|�,U����CzfNM�hN���=$�8�{��rȵ��u?�s�z�����B�rӕ��H{�y�VPљ�洵�32�!FGS[  ��H9Q����	ݙ�i����g9��������@v�l�����J�v{�\f��k�.����,,���ݲK��6��8OЁJR�*����2���b;+ߥ���u���=G�Éҕ��m�����RY	��fj��G�~n�z�:��DY	�@g�T�b������[	㑟�nm�\�8|��ƙ��On�Vf��x�d�c�v�oL�b�J�S� )=n�R<e����.η����1�k�34:��m�;���S�vf������#+���e&)�E���ǲΩ[���0�z4���	|��^�_/=i^1�Xvd��c{=����|���l����腶S���ں�Ku�����N��>uW N]%c���7�6��/IS,�.'-��Â'�� �k��1pI�6UG����vO	
���J}�5��_w꽿�� �6/��;e�5�8��ƿ�K2��"��XU��e]8�:Q�xM��'����jZ�jh��j�&D��K���S���G�SAx+� �kڔ�����c8��õ� ��yk\+�[�(�3����N/g�7����%ܖ%c�Wm'�w)�%�g�Bv0����P)W2�nc��Ґ�]wrDFޓD��҃R�h,�C��g���:��O������i��B�,g�be�ј�ũ��6.3T���׉ �M�%�_����<��+��qJ��zR���y�'?�G���E9~��բ��U�cK����������Z)�=I�p*�EX��P�cojaV��M�*�#cD��&"2퍹?M��Vt�aʭ���4�o=����Խ<��C��&s�Ȣ�5�����j�p*����/�b����g�#Rq։���$o�����6���Z $O�S��:�hy_%%�� �~�B	���XP����Tu�v��V<����LIu�]�e�{k�����;��Z�	������1��R��|x���3_I�1���[j^����6����8�*���-���_�2t��[��z���o�@8g�ž��C�8�RܪSe��RK�r��M�S\���qK4��������MJ=�T�+v|�Mj=�b��~#����� ���Wn��hH�H�ib�B0�G>�ͩ�,1v�����b/���߹������J��/$��S��Ho#�7���ܵ��_(�e1P�c_z���+CZ�m�(SO!�lz�rЮ���d ����<����_�`J���N�0/O/}�T�Dv�h4�;z�>�a�"�\/H����jk�}I�w��Χ) ��v��{�6��4�Ѿ��Ѷ-&U�٭-q��tBv&\��b��Bi=�P��5x�[�F�	Ug�<o|z�b&�9��C�Y��G�q�n�|� 7���6]�El�סw�c�r�ǯ -�L��9q�;Y��۝�;<�}���6���Tn��f�M�)E��1�7
��tk6���:�Qɷ ���^�w�#�*����Wk��qK� C��9L�I�=齾��W��s��(~��ĩ���>�zrL�[V �e�㥒t�	N�gcN k���R�#��Eס\L�R���A�����fkv��\%��3>�8�KwbA�Q{���}���_n~~1�cRP�A$�.��Ս�RbЉ�:&�e�\�\�o�x�X��>���K�JH�!�}��Dj��+��������+�6ޝ�{g�s5&N��s�0cf(���hI��0�v�P��]!����I��U��N�vtU+*��P�R}�W9~7 ���XΤ9Tp=!���*Z�/���:����E��U��k3q������6^=�'Rʥ����iQ��<��f�V[�WZ�N���y<��p�:�u5��s��,wy!�f�Yb(H�!o��"͐]��r.q(W�M���5u��D�;�����ۻ���r.�n:Av/�ĺ�,Y�*-����I?9����m�J/�Gu��+VRm���=Hs�R����S���t�u��U�?��^�af��J�c{��:��8	TC{��C��u���#q�Y�'���g����E�~��_�SsM���C�iB�v��2�$�c	�����V�/<���`f��[��E�l�^�����d��H1�Q��aN��-F�X�hoE:�\�Zw��wc���6���'��ϧsm碃<��'�o�GM>J�>�#c�;�����c��DRH��/~����T.���%���M�v@�R�.O�Ӓ�`��cn����'M�S��ͧxm?f�F���/
�*�=�-ڂ��z�@ϩ$x�O������k��0_��z�����x8Ŝ���z;��R��� ��/;�@s��F^d�2;��:=���ykn�@.F�r �Sٚ����,mx�C7o���әtz�t9dc�%�3&�����)u��|����.�@����ka�#���^��s+�B�mc}�54�.��/7�r*�9܎�Y@��<	J����[7��pt���Euk�=6�:�%���������R��8OC#FP|���vqc�y�?!O�ڪ�@mԭm;#��*�E`��oOW����Rd\�./;�y>���zE��)�{<	�X�"-��n�"M��5�#�@��R5ᠩ�	�[X�&�3�Q�����H��"�Ӓ�I�j���M��~���%d� ����Y�(������ ��>��;Y@��lY���C���g�s{���Ar��H��c���Q�l4r
� �D$��}�]K�yʺI���m|��o��g�����S�������߁R�.��{�rP�]������~�y�������4�ב ��ڊ�l�4َQ�i��P�q�Mx��T��QJ�淇�zƱ��yV�
*W��'�Ķ�p�xy�mf�So��x[�l��������ކP�6�!�-�þ�P�AIP�� ���~�����!#M�џ�T�d�T�T��|�뎫��8%ů<��/��%�F̪�[��f����禔M�X�>�z5j����׍�v?[�����p��}Mp�U��F	��,S����m�Ej;�-G��n����������pD#����o�� |t��]X�D2޴]ІK�����O�4G΅�S���~�H�����+S�føĠ���:�緅d:�$�|�8���H���p"����3ox���%�<�s���Rc�ܞ�Q֯�boq�*�Og@��UM�F��i� ܪ��[��xe���	oW�W��s��x�EF�P���f�	�G�q� ���a�{��&�kc������=���XF��B�>�i�e��?�$?5�S���ތP՞���v��]dN�_l'�^p��c�=Z��\�+�;�6�'A b[Ĵ�,%��3e��+��&����)��؅Y� l���i�>�*#t�@>`�,�ʏs��s����֖�ɍ7^��١��z�F��~ϧ�M1G�!xY����G�D��RrZ0�p؝��KO�ޟ��h�
�.�*��@,ö1��Դs6;tW<@&,W��deeϑ�O�<���B���3\+���Ԟȁ���PQ�$ơ\�
1����"������������[�w� ��_��m6�:W~pW����� >���$�Q���$÷��ͳ���?�`�b�l�ܥ��3�Nnr�-�pt�옐����>��=
���J(�`�"ں�ܶ��v�^�_d*>����)H)���\�||�>?| ��%W��~t*����B�s��N�.��[$�Nﶟ��F{��B=�60�Q����[h�`n�AR=����@KN��	�o�5	���i�PF����S73���G	h����w�{?�zw�$;��������|^6��~g��O��b�o��NP3.$�>U~�i�ݵ@C_���j�
�,��7��y�pр�6���=�����s.4�N�_�]��2ͷF�I7�x��� ���2�M�vK��L$���u�Y��:`7l2��tMw�@�I��\2��}�+S~��N
���ag��y��r�*���tSs�����| �Z��լ��
$�8Ri����n�Cz�6�]�	��/Qg�+gH�mED ���!�5��Ԛ�LĤ5��
q���EJ���%^��	���m !��#����R.!{t�����5�[����j�@Y��K=c0^v�b_@^�_rmOY2�^��8M���g+kT�r���Dt4s$�6d��ں�T���:g��Rca�t7"��yxxL'_�(;���d>t�؞�!3�$�N����Ǟ�x>;�U��o�u`� ���)�L��ǜ>��D�u�W,X�SK7�Q��^6Z���q�j7�9=�)���� N��kϭ�ў2�@�qժ�I)�PSξd4�<���q<����������F?J��p6�PeM��v.3�D����Et�L�;�D-y��9���wd�)���@�+؟�T�{�|�u���[|+j`�oX�Qc��M�Ҙ!p�=����*ǻ	vN����1��?���G��n�neZ� a=�s�â��ׯ�Q."����&j�խ�VNʒq�t����r{���G���O��BE �[���4��k��T�j���௘O��
�;i�'�g�w)ֶ��k"�z+�}}�v�Tk��=������v(����� ���p���*z��z���K� RaB'�5�N��]�\�yr���S�?��$y&�4��v߂�d�Tn���S	�����c��7p�����7�ꅅ1����C��{xߤY-(S���d���O#��J,I���צ���|mƙ���$�Drܙ��������'r�b���t1s�k}�'���F�񌇋�68��
�������.�J7�xQ8����ܳ�F��1Vy�H�߯;z���w8h�Q&9M6�<�]�F����k,�-\��@�A����fk9� z_u"��a�wW��JH��)7Ag���V?I({�������{c]{�n 4�*�l5zZD������%A����Ĭ����Ҏx[@���$� ~I6_���V���d�������߼�ww�$�}:K��4-Ѐ�{s^K����L5��6gv��\(w||X$�}� � �z�OD��GN�я���j����{�#傋}C$T#
��\��aY���g�d�ͥ�)�1����NOt���4���lڻx��vi1�=��HEx������IԖ��؈��cf�70�Q<\hO9�ٻ�c�+�̳��6��N�Ɩ]��<���f!�1�"��/�aPcDo� �j.����e���D�\U���JD����E�\`yH9�L��KA?�NO��C˳��=�u7����ڻa�'��a���m�vª -_���C�\��p�l��}=��g���f���4K�����X2;&�Ű>��6�;�ձ��r�-���{�dP��v�b��SN����ꗟ���Y~�<��9"�0�\���>\���w��;[����S(��fw�r��Y<�,�PUJ~� dS��5�1��G��~|愞��>���o�io`8E�L��;�'�k~�w�=���D(q��K�6?B�׿�Zn��L֦����H�v�U���~���!��;��MB�����L�Н����_����IX�e��e�EuSk�W5�X�s$zt�J�Cl͊���4�e1�?�*���:�+����,�P�a��Y�؀���F���oT<�[�ne_s\���/�,��K�җ����Ir�i�}���^�����O �i�.(Oz�1!�g��>;�o�(-d�l�c����#�A�Q#�����ZO�*�	A�$R��]��l=��&)Ӄ?�4��2/}J���{� ����a��ۼ����i�%D��@�,�t��V#�(a����F�%Եf�)�l
�ߺ��@%{";���N  ��h����(\�
� X�]�ͯ��a�陰��&�!�2�D��x�k�9�5x�^<p�_�]c}f�<�P?�t��a�M���W���o�9�t>�-s��\ S�sw�~YD�	�g�B����)Zm�b�@�2&�X���)�i��w�P���<7�G��̚�۹����7S�k�ͯI
�@d�B���9V�Ց��q�e���2%1VY���c�M��1ͷǚ�7�v�c�+Y(�27�/�����!tA��o��l��짲����'�ާS�lz���X�g�(�=Q�;Q$%�w�e=�i��C��
3�jF�~��0VZm��.�)����ذ�5�ʮ$��,��V��0��JeX�"�u�!-�cV��M��:�����CgV,��ge>�<��i��ߠ=�BG���&��ty��f�xG����̐����I,X��㪛j������H��'��ǥ�>n (�0c(��f���9r�����7Dܖ]�$<-T�q�.D�rT
��opE�l)�(p���m���OW�޹��5��u�<��b��, �����G'ʏ����	:(��<�#�؅�<�	�:�?z�m�>�H���-{�E���e��t�ڟj6Dt�O�\<%�:�������{��������k˳��c�X�vln[`u�6&�Fb�HAI��Xl�ae��s�;����^�h��o������g
o��x��f���АJ�{�%�_����� �?�`ػ�$�[RI`k2֦M���`���gxO��
Z�ez迋����
)-��c���V� �_�g��rœt����hrU��3�pM��徘�~~�U!2*�Aj���H�7>|Si�|Ǹgc�0HI���!�}���OT���Ӳ�t��k:�t*��S�U��ƫr_į_ˮnr������F����n�r��Y�}/|�υtGM(]�?�[���R��SO<j(%b#,�@t!xR�-���Y��'!�7�	�����e���,'��A>yش���6Gb�&)�����{��7wí��[�-�tm����'��j��mU)��e�U�1߸.�"� K��C�z�[����s�'�l��;���}3�)�v�"��,:���Y-j��7@��k�����z�!| իL�KE����,�;�\ɵ@fD� t���VhS��=��i?}}r���:����Dc���%�'�Ye�s%)|K˵�y�iِ��	)'y`��V(Ab����
�"In6vp��,��eRe)�-�I}��'aJ�߿����?�!Ȳ��mS�'�'����~��ڕ"��)�u���yI��q�*fa#wC;e��w�V^NW�.�ɩ
Q;���
k��I'�W��
W���7��D�1��H�Ԍ-^�^l*�>d�*���{JU�@��ڒ����@0%$�İݣ7���ӭf6�����ί逪pt���8��:�-���՟��,�Kܳ�o�sJ{���x��5��GL��h�W*mF)�P r'>G�<�<b�3���v�(�5Ta8��;D�@��6�u�/$�Ig����|��e8�qh�i��Z�M�R4�ip� u�tak�;��Z�i��a�UwFk�&X�b7���I"�Eg�Dq��?}���C�a$�CfeS���v�ҽ��R��w4���������ml�Z�����[�A}�cɝG0����X���_)d������&�(��/�&I���u���<���^ڢ�{7���ZsA�l�]0%���h�8�s�P��X'�m�^�-����Wў�Ȇ͹�B-��A��1;6g��@��%l�d�׀z�@��fX�x��vl�K���,O"r'j�H�����<�~5��pl��S +ſ����w�V���4[ �fe�Ti�}tC1D9���)G������;�e��E�����l�{���L��Ћ��|��50��X�u��]I��K���b�\���_��
�7z��n��;�j,R�����<&C_OA[�I<��A��"MnC��0_�⤻�و�ޮAZ=��$%�N����19���ؓ	�ՋwW1�����UH�V�I��m��r\X_uI(��?����+)��*�d�壙�$!.zNذ����N=�ǫh�V��ϷR�������k@���!�jG��K* ���u�߾�$AX��K����f��ϔq�B/�p�ёE������WdK������	^`-8:���xl��K����*��ɔ'8�:!�������7�!_�v���v�'=���F���<w-;F�p.Et����[�����L-�%�''���7Ypv/�'VU6&���wR�!�)M�7��Y/��r��Z�V�\�_�~��?��q�?���(s�sn`|�$��6U�JX�z�H"7e�_�б��5�e��Ӛ�D��;	����]s���G���!�a�P�������f߂%�j|6�j�^p��%��R5�S�b����h9�j}����Ȑ����p��(g�Ō���̼�ю�g���E�ƶ���<�&͆���һq`4q�Mf��,yBt�a��+m�ڶ@�cў�i�iX�h�$�v�3G?���<A����e���'�Z�Z����F�ō��g��`f�s?
��]�� |�6��x�]��a�ҟ�����}���z����I=ˬ �չa��Y��D��*t'L�?>�棎���=I���	N_\~ݘ����v4�eSoHqDZ���y�z���PDU���5t{��>H�\*1����z�	�*"_�����L�!�����>��~��eô�pȦn\�֎)������,5�R����}�>��kI��kt�BV�ɫ9���1�;���@gvh@\�=��(��~��I���rOOʿ�����կ���߿��]�6����C��mY����������5�d&�X1ӄ�'����⥵����ݏϤ�[HNu��ѫu�!�����M�*���"�Fv&��������8><�/5�-l�[�m�x��c���!�g=0  (�*<��X�0`�(%�����(��r��w�xq����|�v�<o�J{�;�A:�/�ܧX�����Tf�1�����U-�� ɛ'ɋ4ck��q���������,�L���Uz�u�PVN�k�<���/+:D��ߦc�Ñ��Z��lO�4�`w++(�rzY@@ to��
Ao�<��%����>
إi�3WK�'�O`���I'���5�a�n��̥�I���7�ă���ݝM���i��+����SЩ�9��ϰS1֥�_����3Ks�*,��e��h�Kk�6'88�� �e�`���NVz�=f��������G����<���?u5�	���,,T�;�N���{U�R67�����6��A )�E��ޘ?�J$E�nZ?)C�e��8�&3�U��E
/��Kr��K��S�U�Kz3�Gi��o������&�/E8<=�b��:8O崹q�UW��`�o���}q�'ؙ+3�����M���ރ��߸ͭ��S�S���~��u.��.�R��k��H�)�륚��G��T��lݘn��[��<��l��+�*��3���=ϸ���g�O�GVH�6�9���C���`���?�p��x�rJh�|���S�h�aW~��.X�)4!���7���1�=�7��c�mG+xe�lڍ��伴gnE�K)�[��rV+�#x���T�\��'m��ڜ<ɕ���ѱ��X��Pӭ��Ŕ{9��H-+����5�m�ޖ��/}�Qqϒ9ޚU_���t̃WOZ���$C�g�_����ض�)�X+��(~� ʃ���)P�?r�$��_�$�|b}�-�Q� �nҀ��`[�nҚ5Β*�`sz6��`{w��{�e�|�(� 2Ra�V�^~0�3�xkM"|���g�,jH�`K�#��g�,�%�=���#���_�&>�A��O��RS&�N�1]�h�6]�zٱ��v�{��D�f1��ef���ᚚ��܂f�F8�>�6���cp ^p*��0jedݖɋ�y=~*��:E��'!#R��}�YҾK}�x}9W��,��'�S�q,�������wwvpڪj��.��~~�M+���*�V��J�����X����1�_�Jg��#�P�S�D"NPWBϸ{��&I9'}N�Z�_��DN�����=۹75�E��X�E	�ã��o��M��/	w+���Oz8��X��'nw_�,?T4����@ҳ��%^`��@���-������V�����#eecf}���l�9��t��T����x��	�Ϥty��$77��F�[����Ҷ�2����[�⇗:�~o6N���$.]ힱ�t��&� ��v�񙛝��M�!9���AU��Wh(�~U:`�)w?���A����K(�"����F�+�	;�9ztfV�k� ���֚9"}�	=NRH�����V'�C'���)�����r!��{\�d�t]��g�|Ɖ�,���sU��j|������M�)N�\S�hXKW$���C�(ljk=��u�I7vxl��@���qi�<��%�������2U"
���03�A*��'�r)y��n�yV$g�0��gF�&��)*vmo�4�(N�����D4�i6F�=��|)�ȷ=�̄��]nأ��T��y4�o������o��g������56LY��z�3��'��\>p�"e���������yR����u�H�ǲ�P�1�����`�Y���o�|X��I.�,�5��O����/s��P\0�F(��D��^dqdw�,&D�z�`��C��� �h���q��~m��hO�BS��C���]g����,�45$���jғ&/E��s<}^M|	^�l�RZ�5ڭ�;Bw�$��	�޿�(�X���iNi��,�D��TN�!��8�#p�]�Ǫ�'�J�.t�&��]� 4:ofB<@���rȪ�����ϖ���6��A�Ӭ��0��Y�#q#���K�����x�s���w��~cc���@�+ �N[�vͦ���.u�9�ۘ{Hm��xH���(��v!�I<��!�"ծyRS��
2Ƚ���.@+�䂍@�d_d�P��t��
�M��-���Hq��Sخ�5f��@�Z<ՏWK�+G:k�ع���f�^�%va�J���$��9�Wᣱc��J��
a�p�)��/H�M�΢��|���X�X R�����՞ڗ6���Z`�G`�%���� 﫥D�OF�þ��k�}C�Pg휳}���w�<��� �RϾB~���J�pF�lM�z��w�^���9y7�u�D~g�J$S�EH&;�z�K}�6p�k&UD��Kb[c,t�/�~6�
��3�_�w���<">��0�[}���x���N�E��b/�����$ih��O��>���ϖ�����u�ik�%��߬nm�8�������p��NL�݈ryY��p�	�`-��{��HQ�C���y@Cx@n<���<�	ߗ|�@:/�D>�M+��C7����#����qH��A�3���z�>�����SV�����_��M�|�gr�Y8�iD�f<��p���@�D��ט�\e������썴]UX��|d�-D�p%b"X����k��D�������Rɪ���t�N}�����u�������V�x��u�n]5�|Yp�VF�8�܏'L��F������i�<>>�}-3���<��&��歧kN�Jwױ�2f�GSC�xJ��� �K�
���|M�lT>r���]�>�S�ߊO�J����w\A2c"�`��	�R3R}���f���`��UY���+��("N�W)��?_�*��
VK��֤
�5��[��\R;u��%=�q����ɹ2]Պ�q�F?Deܻ���מ.��ollB���w��G-^>Eʰ�8����H��t��{s$^������v�*���r��F��o�E�6��b;���$sڷ�sD��cߟ�bV�	��~_[�?��;'���ˑ�?��#ۥH��i}�[�`!���g�B	;r�TsF����`/'dff�~�IN�o�C9�ݱ�l��[-W0�WhO9ŕ)��_%�zqmm��t�y�n�R+x���#-8��u�N�V���D>qS8U�˒0�2�ɥѵ��4�/��[�l���NIc��$d�V������im!UUݕ�N��m��7��^H�]8����[U&�k�`�3���I�Pơ�0-���L2�nVœ�b��Α�O#�
(�nƶ*7m�#�O .���8݅�(��ڎ�VJ���U	����`kF�؃;oi bV�ɘ��{��+p�z_���"f��fi��h��\����yQq:�/uU���p���.Q�D���LW��J����,��_��U��E|$*��
���&��v�� l_��݄�FI	���v	��m�gW�8�� 5�q)�B�����bDMG�S���e`��t���ڍA�|3���������G�y�|��\.w��*ɮ~N��w���R}��}��A�W���\^������@��*�η �a8�������m(�\�;�d�nǑ�vaF�R�n�O�Z����h�M&d7C����ɓ��~aa�YY�i��p:.�3�S�D
q���6P��s�K��S���_�E+�Z����`e�/�/����!�yQ5��5�T\�A�撩4*��>%zIY�SUJO�����������%%%�R��t����T�M����"s��O>G�������."�t#]���HJ����K����(JJ	K/�t
H��.%)�t/���������Ν��<�ܹ���m��+ݜ�U*��ӤU�4��>/!d7���,s=������N=����D��s���%C��͏��P�CS��F��$!pw��N芧r���[+��������Y�v����D��[9����\�A�dmmWe����>����|��s��y�'��<�tg�y���N]��;ő'A��#��њ	�� �N�w�(%���(���TJ^S�����m��$ţ�ǔ��U#i���+�<{cs��r� żK� ��@�C����#V��E��i�F_�|���h�vF�}f�m/��L�~���%����<_��ff��g��9oծ������(� ���2���D`�CP	UR�)����kǴ���f�<� .�K���(3$nB#4 ��?9Ҕ �Y�<3^X_YK͓>�"A
��9x��M+ �%'�Ɉ��=k���ѐ��8G�6��q���m(Y�o
�a�� ����62:�M��xՆ�t{hӝ<"~�g�m��%��fXy
q�X�����lz��O�?��!�x)7h+�u*c:6�����SuU�'�#���;R�o���A�G� ��?t��H��6H9��ʳ�Wҭna����<�?��7J(.�կ�o���J :5~��?�Imy�˹q���.*!�Q$�������U�"la�;����a�u����͆RI����}5933��'��X����zza�W��-#M~���60d����2a�ZfO��5��W�?eWQ�dP��~�Ϩ���;9 I���QOn�H�G���w��z3�=���)������u2���'hUm���v;�-ak�����ηtg��aDћ��Br���k)��̵Y+Ƽ��,f���<u�$�'�,g� ��_t�اII#�]�xj���]��ah�t��A�%W�I�,�4 e�rU�Ҳr҅�V{O (Y8x��YrETP�3��2���q-�,|���W�`}ǧOҽܸ^
��D�ԩ�O��)&2�D|�p���?m�����⽹P��ĽO�=�8jc�?�
}��ocE:ٹ���G�ăc��ui;�ރ�#�k���Ԩ>�Շ��d��&�#�v�ф���|S{3�0��_�i����qEk���8�7=�$�ɕ� ��~�lb��q���$���ؘ�bE�B�Gd$2A��t�vw��*B�æWUQ;=��QaeWi�r��f��*�-P�C�v ��ƾ���6+y�=�b�hSr�-��T_q�_��squ����Q/d���A���K:ܮ Gr�N�7���X���]�{����6v�� ���v:���0��+S7�J��1�ʻ>Z��FrK�*z�|��8����_'ߗ5�w�"kt�aMlC��O��d��mxi>L��&B��Њ��?Z��C��=�� v�߻ᡷ-�~y�f�X�:k.^Iى���sI�G]�n���XG)�Zz��'���;NN�aE�'���}@x�D����"9(��(qp� D����4E�|K���bW������|�0.k.�Y~��^B�H��~�<�¨|�(H���ɣ��7�/��Ytէ*s̟�O��xƺ��+=�`33�A�י��|��6w��!�H��d}X%bz�]ߠ)9+aO�&]�
Ĉ��+�%^�����r��gB��&S
?l���S<~���[�^�?�@�d�|TPƜ�����4| ��*�!�s좭&D�U�����e	f�w
ǥ΍h.��4ުCުH�}%�妡R'���^z���.��	�_�I����D�z#���r�E7�W���{�)�\ �����3��R#9Vq���d`��B��|@�d�����AP߿�v?���IU�7Ӣ�h+��������3�Sv�F(w��y�f
��eh�kF�;��{��J�,_ҹ����%� ��&hfN)9������2E紧�*�ԃ��KJ����������HK���E9���O+�:i�wF	,M��$@P�f u�L��Z
;s����7�(�d�Y��y��a+�4�b����_��	P�a��~maى���Uf�=RaQK����U;GY�d����w��uH@ǉ�v�]��CY�T��-��4|�K�x��^1���۵�=�����WM�$��.M'(��I�U�����yyv�@��=�<M/�aPnq}�3�����Ig�}��ϟ�6���ĵ��{����;��J�����	��q,Z���+
3���h��i�ӺP�=��gl�*i��8x8Ƕ �����z&����H���Ŷ��b��TBDz��a�L����Ǚ
���k��x>�\�z.<������F[�,��Ǝ������b�YCw�V���c�������t��jE:�L�y�\U�?*r
x$Ɵz:%1c��:g?��>����=-�'���$tD��E��I�GO�$<��� �����p�2�"�Pܶ�X����p��/��m�_�����{�a2����Ј��?i��,�P���]�^`���ͫkj��-l%YDBL�k�YN����O���Ɏ����:dV�1��'C�#嘉M*�:�xc�Fۘ���04�2�"�M�iRۗ��'�]��|\ҟ�di�7�Ѹ��jt)�O���̢K�A��5�0��qҰ�Sp~k���/�<q���?���"bg���u�P�yWq��s!������o=&;�]`��J UB���^�O 6����Ğ���Eu����}����U��|������L+MM�i������ע�F��̃�[g���ʗ=�ҘWnKz@����s�RvK崽�'=�h�h7�~��������������qE`V���+�O!AS����A��q�".�����_r��<=�c0drSS��\T�F}'�-4�2�n�;�S�$��N7__Q�l�{����>���˦��*��]H����|�z��L�~Dr��X��̚8PB#�ý�s�A���0�|��+D� �L�3A�5���g��5�}aa�k� ����,/N���NY��J��+)V��6�!�;^��7�L�pXe��E�ǲtX��q�t|o�~�jH�V��"S���M�#R�C������v�V_����!�5���i"�$�瑀ω�1~�l��U�~�qC����B��x?%��٤	4�z����+׻/V�W.�S����g��{k�@J��ʠdg���ɐ��J;��pq�����|���m�т>@zk��e.ψrB˳ ��^V��	��� w�5yrR^(���	�����.���q,��������zl�̽�TE*47�|q��N|Ez��y����m)��e�k�X����R�>�91
�i[���ߜHqw0,�֧�|:����ߟ�<���B]���7�jb��S�I��-���R�8�k%O�;�6�=*�$y,IIh�4
� 8�*��K��r:3��(y��(�LF�F�����S����f�`�_�f�6�]���0�(��0(�??���a6�28��b}1��"��c�X�"�Ƣ9�x����V����n1]f��ͅ�Q1���7U��9�?�f]I��!^�E��^���D��e �����\�2^���	�	~@T��.�4��v�3I0Q�7�ka����0n�����9y��������q�ύr�B���+�Y仓�(F>+����zXbzdjj�	��L�*	����!X�G�/# w�K嗦H�����=@������:׿�V��l3T�e&��8J��:M����]}�I�Q�ۚ.Rbv�P�"_a��[z�lk	�i��|�$�%�R�{����[���Ӌ0�N�v�0�Q+�U#��l�*66v�ތ�V��fo��o'�]@���W9�K�R�����T��hN����>͡���U�w:��2�S���2�� =���Gl����R8�Ks�9����a��EQ��'�z��nP�7���]����+���e��~J����~��	+��@X*���b��̌j�#P��[��)rξY��L�˒py{�C����U�i)����5LZ�ꬋ��`^����M�=C�����ќS����2�/p�,�]�8��s>���i�k �2c�@R�oR��#s�����U�E�S�{�o�]�1c���
H�_��+�<��/�v�N#A��a�	��'���Rv��1�A��'�޺���]N�ԙ��U�t]|��� �NL�Tץ����������{�LE�j~��`F��7WL�	:Ó�X$����"[ת�k%)4�P���P9T���@��a4��OV��vi�Lu|;����t �?��պ��*c�d����~��܈���i= ����0A8�{�+ŻK���baqr0SA	�E�>O�?�:����%���o��_��) ��97U�D�T��!�������S.����W!�,,AA-���a��ʡ���-�s�����L�y�~	����5jS
��N�od��kMh�</�I��*Kj�Fk(�=�׫_2s~�|$�'��!�euZ����D@�=���;�� ?v���~Dnf���i9cy[ Y��239r�f�zv/��[�1��݁_�E��e��8
�
��K�7� �ER%q�"��}���Jo�nE�*�n����P���o$[�/�s�붖Fz��5�҂���r%kٔ���^U���h��v�$���{�/8��yl����KD��E&x�0c�بa���T64��W�P����8�L���A�ǫ����O!c6�O8 =���KO�Q�~��VwT��kw�;�m��	�N0c�z�Q>3E�p=@�u�#�f�}[ΰ������I�N���c@�)i%9��rty^�4��K@���V)��cwW��~��+ϻ��~�кO`��i����c�Ba5�O�"�����z绋��N���6B����jT�fNg8�W��[�k�A�W�߃C��8��"���c�l��F7{�X��I(�3�x����]Z���Y�Ã;L��2�@P
�5;�HM<�����x7�;y�9�c)��j�
�X?WQ86t.��\�~�~ �e Iw�P/zIpx�w�D������2������ȼZ3�#�+Dj�-���Q�D���ŭ�`_8�ց�%w_��'�>�`I���""Z��YP�e��췾'�=�ߣ�{�����07�yF�K�9������	E�Ng�Ӻ���^R���B�tk����7���Ӗ?5�7b<6�!���)Х��fu-gV���!�3�1�}�D9��PX�V'C&4@�O�V�D=
�r���a�S�a�X�V�$�ٜ��|�Za&�MJ��잼�~�?��M�\�~V��''i6�ٍ֭��Z�4���D����I�
�K�S0�S�S�%��Yxy�V�"+5�����&�I׻��쾂LjOAb})�y��q��>��C�Ahs_ޤR���}'�u��t�n�����@�7~$_��G��NF%��;�T}3_AW=�6��OW�L����z����R��}[����P��G}��'�޳W�y\s:��I�IO;7��4}'��᳾�7|�W؆�VR�e{1��Jw&�9W@#C���H��G� ����tjJ����c�֔��Ov�p���fn����T�=9����Z��R�`\/��y\�wH}�j?���U�N��%�@�y)���C6����w�T�\#+J�m�ɽ�K
4�������
�N��~�b'�ؿ3��M:� k=�Fퟔ2�[��J8�U`��k��o[]����Qv�z��vmhh��z��_�)Qh�: �����!IlL����߇�o��J��_1L8
��J��ޫL�̣�p�bX�s|a��Tq��AՎ���{��l,���ߧ��zi�W��''�PC���C����
ܭ��x!���o��s׳���?H�7{p;KCތ�RU�iKL�N�yw&!3h�d��%^MC� �?{#�֣L�y��t\����I�ҵ4�>�pQH���H���9�|�N� u�V#��Z�R~pdW�l���E'���������?�����F�=���hV-��I�X{�Ի�67��D�b�cV�\3&�+��~����>�ݙm-��q�]����a�I��x�576R����]~�/����CH��x2�~3 �	
��rv�e��|#U~���,��H��r|�>�@�#������++*,n�TG1��n�77�������
�ٖP\\�u��HK�,����Z'346�K��{P�T�C�N��;/.���3��Z׊���s�-�M�훭��r� �!�rd�0�ef��I\��]pӒ�b �n��#ŒGY���fN3S䍶�|��\�[{���c����
�~=O�������+N>��\,xdu��Z�Q�R��4���~��� �O9H6�+��?['i�3��Q"&Ǥ���z3H�cI	/�����3,�B�E��FH���tI�޶d���,A3S��.�T�/�e���x���UQ�ˉ�ç����ퟥ�9�~O�� �PYWgW������G���K�����o�������nN��}�1���Yh0�z�5�r^"x�9xy)�U:��S�uo!��S���C 姫'N�6N����Y��@uuV:�uR~(������X�����H&Y�_U�����o��"I�S��u�������4>�U�4ޔOv�N����9��1��[__oPs�tJ����m�t5(8�X$�g��9&>9'��K�!d^/��2��05��xX.���s9[������9��z����W�K��qo��c?��=���N8�������`�\ӁM�����rv���]���U�{ɪ���eѩ�0�A���E݌ȣ3�!�s��5o�W��-�P�^�1ˆW��� �wSk��h �h33���,my)�jSUE�cnBf�%aJϺX�����?>[�-6��y�j��q�$%5u���up��"��
d2��u*��1\�,��I��v�X���4�N���J��L��,L\:���t�O��m��-�_����,	;���R��F�u����kà(���iW��v���]����5܂Q�{;54�8\O��fw� \�U���듛��K���e�����_�������egd���p��*���,��I~_��y���ȸx�B�_`���}|0�0�l�F���<t� _�� ߢ��ak���!��n��u���S�g����LO��]W<ovM�H���W���x)gn�U]]m��Է��i�e�\�>�A��F��O��=�h�?Z-8|�}Ju����Vl.���V�C����.w1���5�>�;LF~�)i�_F�sٛ�3=}�r_:Y�Ԇ���who�>0���\Lpq��y��q��{�b	6�7� ]9���q���	*�~���+!�ĻS�j�Rm��ǘ�"��Y�D��r_�+P��X޸�?0_avј 4�0��������wB�>�݋���ܤ�̵����R�w%�픈�봪pH�;P"J����k~�Yq�M�f�h���"�i�JM�V�e$Hօ5Id��#@�]Igu�)@�n$:Z����㐬0ˁ��Q]�̂����U~��-َ�$J떿.VVO��7�1<j0��~�����-��Vr6�!�a�S��i/�~�5c�4f�/al,���"��⽼�	���j:�j�kT3���M�Mr*��<؊}f1��<$�U�~���jໍ��+s��8b��aW�E�V�6�6��u�R�=?2�x��M����C
�Emu�ѧ_���=%��3.ӯl�Y�l��B��4�ÄOH�Ŭ�u��[Qxs�*�XF�����I,<������,7ifO��T1�=N��F\�s�Ie��-,�����^�qz�	��䋪oP`��OSÑ�3�F�����&�dP��](KF�(���m�cg`ȹd8�v|�`:�7������q���^n�D���@rK!��>�8Y�ڥ8���7��q6r���Z��w9�������z~D"�h^ب�uʎ��ˍ�F}�_T���%3W5��>�q�Lv��
��7� �����ͺ�(��،���#QO)�!_��Fo��/ˮpN���z�Y�F��9d�_�����ir5�"�L*�}�!����bɨq�*WV�s���?0�]�N>2� s
�2�S�6�mM]��ߚ�:3s�'��	lD��S&v����Zf�P=���1�ۡ0�+u�ό�����r�;�˙t�ΣA�3#^Ϗ��OF����
����~
�N���I��D���`�?��	&p�H~	���}A���q�[�b��:y�.U�6���'
x���ׅ�~,��2+�h�@����XV�
�����y�% (}wqʁ����,IU�QH&��UDЯ��웤��Mp����(��X���o��(]]wث����⫊��(�R���G��>��a���i
��b�����o��2�Scs3��%>���<FBL�$�}�<6�ۛ)�����_+�$��h�JL�+mD5���w?Cw�lW.�F4mL}Q�?�~�8�>E9�G��6���(	9?cH|>��M�v�@�MAِSKuI��މ���c� A�T6��	���<weSv�/���Փ'�� �^��4��mZ��5#-�h�tP�-��o�ow`����ԄW�ⷢ߮z�W[��tX��$����vǫV��MLlz���n�F���V���R������Jl���h�d���[v�/u��o�i�]zV��K�@�̄	H�~�NX#cEA�ew~ff��kYk_`q��R�/�|�-<,��/P�EAi�Sp/�7uE�50�T9��M/�M5j!��R����bfH�Qc��pH��i(7e�!�� &S��˨hu��:B�qH[�0M�BYO��R��m�ST1�ԯ��HI�޸�ΐ+A'��O��	J\)�����`:���a�H�Ϋ���{�v���1'����s��a�8/nK,�{=/@��`�4f!����c��M�Y�"D�n�<vs�?8�?Ľ��� X�DM3�مE�39ʒA�_�vM���AU)_j�OX� nIE?�*'���������)ۈ�����y�ۍ��Fl��0-)z�cM��?�L����6q~A	K���W$'�A��T�լ;a6�N�s�[tV����xL���4��E�!��Sl<1��gݨ3��k���а��03z�q�D�̅��7��ք8}0�&:\�Y�eF,S:~������x&QrV7�.��zq�����ܬ(�eA>�"��#͐>�T#�i�HB5u#4�,�n�V�u�6�:�����/p���z�t!4#rG_����!�ɂ�~��z-�u��"� ~�a���r�/�Y�؀p�WElU:K��NھbR R�C,M���6`���<ڝ���j4D9�xjM���y��t�8�+!�l�m��5?�[�|�K��:�}����vzJ�����"fØ�F
��ϽI~ҳ)���y��b���3��0{�Y�WލT%�^�~%���m�����3{��H?�½� M�uN�!<Is�#7��JE! �(1�#奓@|�UݏN���k�'!�]�c�_��DQ<��<S[�|���d��Ӆz�j��J�C��$3Q��r�=���}�w_�EQ�}Ѡa��#��ݯ%//I0{�oH�����q
�v�:�?�t�"`����
௼��F�c9O���/���܃v0�h��x� ���j�]y34 �ϥ�α{	\V���SH�;!>#�,�N�|f�`Ԇ���8���^Պ��/�Y h�v��j+_T@��W)�
GuاoiL�?VCRA����G8x5�ix���M5��l���sNz���
~����>WN�-s.*f\vK���Ɠ�u���%%���b`+�o�- ��]HS�`d~��W����T���D��)el�h�gz��׽癛�?4�M:z{f����4�F���	}}�'�06��v�|��ڍ���z�N���F��^��*�a�mt&�S<�V 12��<�S�/�
}`��AF�8�35=@��b��P�H���
��O�dh"9A� ��hz���^�pE�#=P7I�٭�Yn9g��E	M�7�D���?��4��V-\�}�dH���_�=�
��l/A��|1�/����Î�i&P'�/�t�^��]:fw��^~�b:;���k����9�k�/�� �����^0tZ^����� "�#��i{�[��;���]J6J��O�(E�E���L�͏��Z5}���R�
Oo����l��p���i[y���I�c`�;��Q=$ƥN����ԛBPqbCK温�ow�H=@�zn�ޮ֨#�hs��@jx&IB&=�3�a�����}�X�*��ԭ�QRRo��C�t0���~�l%D���!9f�9�Z�3��a��w��2�nÈs?��)sw�:;-�Ћʉ�����y��v-��O����^����Qra��hhX��׳)���=r2��3V9�~��Ǟk�& �u!N���פ����I�MB��Lx�Wg����Y^��m�z|=G����n���(*��x����M 5��k��� _N�
���u���A��!PX��q� [���b�'٣��a��T9s��׍��9no:H��c'Γ�RFْ�l�����}���Ix��,������%a��ӯ�E;�hZ"���r��8ā`�I�tjv�����mI��
㲷>9�^V�]��SoY�.b.��Yj���l��>p0�>󇉀�)2���(��ӻ���^k�鱃Mj���d��� ���2���?�Ӷ�����Vr�{�C���;q�����g�9�;�_#�g�+KR�[�W�?�Y�����6"�$�Bd�Z�*�Ӭ~��@mo
��؄�֊��X���b���_����Y`B<�ă��FW�j����ꄸ1�)��̸kޱ��V��������h�}b�i,�5<O`�t{���ʐ당|�ԉ���)�i�\Y�Y�����]y����{���(�&�S��9���va��ڝ��x��	KKr���2�=�K�>�v���2T'��� 4G���T?�F��)�zq�M���VE��$�e�
F�_e�rUmi>��~o�pѩ2�$���A-�qߔ]Y)`a�/��L��'>��K�E��Ta�O��P��E!�2��'"y!@���L_��'���y(���'}����;9����؟�/;=���͵�e������8�B�`t�R
�wM�Z?[�U�v��W(�����F�W����@i��!��ay�[�����0=W��q�e\J���d�ȸ�a���WAo�q���G{g��R\c[�M^�>��@o�<�I<1^�`�ɺE:��n�����H�+��cE��֌w�ý��-Wq����V���{%3o�_�P+ao�����ݴQ1?r5$vss}~6�I������bo�z�G����q���_șJWJ�3����ย�GDj��BmS���+@�Q9l�KQ/"ԍ�.�ՙU8���b�5D� ^�"��w�1,���[{5��?VkC�n�Ţ�#��O���7������F�C���}U�҂�E1QM̽ny���C�l���O���%]�8�|��JW�ٹp��E�7������=���.^���my��=N��UQ�B�lTߖ��KcR�Xw�p1ԣ�A��.Ja����pzo#��i�&K��`d ���媟l�gGϭz`F��-�vwZ��b�_�'��k���5��'�fsw�2
�`-�w@��e�ט�$� ��͇��ݷ*J�Q4��l/܀�5ݛ�U�>�����z���t�������(��?�u�;"e	��qj���7(vS)�.��ʶ��:u�9�A%5S�P�bQo���ׁ������D`I�EupK�6���2���4�Jg[�l���*�Q�$������Z�ZiB*�r�91�iq7b�u0<�<�f2u�"uڱ�G;c0J�)hv�MGǙ�x(u�k�o�"mo�b{���n�!��L�gV�]��{A����(�~��p�K�}����S'�*B��4l���>G��.Ԇ�˷�k�E�t���m?m���E5?�S�e��S�[��_]	}y}�e_�jPgG�;����ț9�e]�N�3�'XI��@��Z��(U��Z37���SP6�DJ�8�\V��"=�$!D�CNL0.k��cO��툐?X�ϬCsJ�a���/#�E��݄l�l��vq��򉱘-zl;�LŪM�M�6׻��J�ڂ#��7��>�	V�p��-u��.�J O;p��k����ٛfx-�2o`s���n ^��ڹZ�ǯӀ�^eҕc��73����ڷ�J��r��2ɟ�|�J��?˙�Dg%��KWא���f��dG��3w:��*j,��r2i�E����]P�m�L���$�)KP&f���
@F�^��6CR���L�b�u��l�&|ѱ�V�� x{
"9D^��fG"d=�?�"w�a�&�G�%����Z��.]��mp���O^��=��Q �8��<�uN�؀}�2 l�+f#�m�:�ރ����J��3�2?IY��M�
���ne�/e�!˾ŝ�.84@aw� ������PVM����kO��^�/<d�N�5s�9N����e��O4�Dʹ���C�&�[y�D�@�[�(U3d�	)- ���wgb�A"����Л�o%�����>"������C5��]�N��b���ŇL����:(r�����%+j�,����SH-��_q�g����G�����m\�ƒ�H�tV:�5E���CP��X��c}��ƺQ�UyiA��an�ū#��+��R����u]* �{�: ��3cv2����bTء/�&�<�"�/eP#é	��+��UM2 �a�&�5�vb@�p�]�dB��MZ�)P��������2(��8���'E���T!['���f�ɪ'@I�X8`�{���@�t��A���[ǣ���o�9�	���f����X5�9�/f,/����]����f�J��Q|c ~��۰#< 6�pF�ӂۡ�I&r���ȇo�zxx�DL�Ɓ����*n�@�d/� (��5$��q�b��S����̤s�#�䝁�,��u�K��MB���-g����r�M���6�ۓM�p����7�S�hܦ��i�����g�1iN�fH���~�/�����LlaQ��L�.b n��B��i�UZ�0�i�_��~�V$�q��H]������EIxD\VXԣ����OJ���ǃu���dE"|�?wށ��[ZϢoR�����ֳs�i�7t7�	�-o48%�u����n�YH"�k�Gks7�6�~�)�� �jR���/�FP��ԓ�,��I���c��csĩߎ,}lo�yys�4s����4z��\tw��l>��6���+s{����$����A���!��ɱ���ܤ���9��zUX3�q�.�����_���n����o���2��S�Z-�L��,�%w�:+���O��S��BXi�;�����d2�P���t��X�R4��L�Q�/dL*�.[+�د׉k����n���g��&\ ��Z��-f,Mcv*��u9�l,ǩ"a �x���,��o���Lihii�|}�
�T�C��+U��RC�6d[���\GK� ����1+�f,wsiqY�[����	& �+l�
<�"-��9.b[m��[\��^m��lP�5v�$��;��'������U���M�����	-gK�W?U}�7��Z����BSO�Oa~�^���_�%�W
�[/���w
@���A�;l������>����6�y���S2�Ѽ5�Uv���ԓV���bh]7.Э3Ίy�?7�'��c��O��K:L�7;���,���� ( G��bo<����u~Ŀ�;����Ŋq{e�͙Ok~��avO�BK��yuKy���IɎu�s���A��Ϫ�G(��vC�f��#��a��L�^'�\p]	q�yk�����rצ��W=��s$W�jM�Rsӆ/��q�W����_�g���Gm��Ϗ�Zm�r3Œ�O�g������@���E�e� ����C�T5AT�"��@j�;�rx�qY� [�L��P��+00��u޷���-YdksKNj����,Utu_�>q|� 6��;Ώ�B��|yjFo+��*PR��o���82Nca�%���sF_�G:��#����rc,^��v��r���Q`�s�������]Di�����l��YV^A�#�����[�_-k1�@�{3��������(���;�ަ:}G���A���<ۅ*�N���~�D�+P�1@��o!�o�P�S�!��f��ld`R����ϛc�wv��]�5j����=�����E>r��b�&t֏�9i�[�>3_EQ�7_��46��ޫ��I\��F�Uߜe/����A��7���k�V�����S�Q��DkCC+���9�֫���`��������:����	����� ��5�����ǷA'�}�^�|{6��=�8D����d�,�ۣ��.::�����ͧf��c��v|糭�s�Yǝ��2�jtB�l���1Qr@s�]��'��焪�VA�ˤ��*N��A�r����hu�q�­s���EG6fj�꓏=c���n^CP�8��sٔS�����Y�;or?@k���@eOA��e}�'A��o���	���?����A��M���Q���-�2�m1]�n��Q���w�Z|u������͑�H;K��_��{�-8�J���Л��sް��wD)�!��'yo��Zi���
T�}�&����K2��.�܇����p���эq���������a�K�)un=5�Q}Ae�}p(�)ߘ�zĸ�Ɲ���UY�Y��T�5�C������8k��ě,�B	W_����=�����1^�~�U?�(�c{���7�:�L-~TGw��R��u���I����+#��d�T c6wa�e� A!vD���{@3����At�����ʟ����~�ũ�=ٓ!oU�ۛ�>�@�A��^��~���)u���O[N�8>@�6F��҃jbﵲ�������X����'�N>�X�����0�c���,���wCtV9��7��4j�v �_|Y}-tn����n*������v큸����V1a����G>v}�2bZ�G}�?˿����Ϯ�������0�N+�&Ű��҉*t}V���~�O3�Ker�����'@|=��V�矞��kL={O�Gh��%SdT׵�N>�yB	�0�`�v�����m�T��8�DԚm����S�_887���MU����F�o��!q���Zn�aN�e�@w8��[ҿ�����Y����R¨���vBo�%���yW D�!� �eQ*	�gi�Y��9���l��T��I�>O��EA��)��U����^��7�C����#[ǘ�Ҕ��{e��,`��rL�����t���Y�!"+�ɱ�� ���ڹMQL�B�k^�߁����5)T@`��n�8�'�7hZ�&�J��l����Lwd����r�H�{E⢽7���.�&s��K�;��폤A��=M�� r��H���Jhe^:���s}�A���J��e>M�I��E�P�^��gs���O���qv�`ߝ{��8�^5��z�@�D����nM��R�����z9��^�8�;�+��NǶ�)�2 ��5{Sk��9Tv��sӶ�=��[�B������nW�$��;�x��=�#8�Ы}����@�|�v7AVs̮W���C)�}�ؠ�����#���n����4r��$$�இ���?�k�R���A0/4Ͳ4�6E:� 9�p�fS����_z[母�&�;���R>>�ݱ�'�'j���6�E2���,o���H�Ɵ�O~;F\�_8��3|�8���^�`����ǽ����P�K#6'�r�7����a��а����o(���Rvo�w�02���Ĕ�2}7m�2����i�1b�qT�N�EO��{�gS9_���N�BdM~D�c�E��9��O�F���@|8X��>`j��k��jP�����+���a4n i& �4&�rs�z޳��̱\մ��>�ϱw�������wCYC%�����B��5�-�k�n���0T�ԥ��v ��}���I�߽���NR�M�k
�g�����:���t�X� E���^7'�r�L�f���8�{��wH�Y�q�P��mw߸�C��z[�ȿ�x���/%�Ma�CP���m`T���ז��1�O�A��/!������ 2���q����ivM�t~-%���#���i+�T���\ӿ{�a��kx��lnݐ�c�Q��n��q��ފ�_��b�,�L@B�F<8("�x��P��|,��}���ا���������`�M�IY��,��DN�X��4��E��.����*6sA�x�n�w�B��^��t���	�鬡ʲr�l��C^��*����ܜs;���l|@>���W7b�.�,l.����ZB5�p�z3x�ov���V�jZ��\�Z�<���ޖ�`�O�3�f��A���ֆ�f/�9��j��4��hNLv�$},���-����=��ٜ��k�Ǣ���L�tu�b��ih��ʷ��_���.Ao�%�*[�"Pe�+H��rߺ����U}�!�PO����Z�sV=���q���z��T*�L�Hk�%��hV����~g�.�����Y��L}uT����"�H
()R�A7̠��tw�tJw(J=)�� � �5��м3������`��9w�}�>����}�T2j͡Wf�\X����v2����1v:˥��y��F��\��䢒��#Th�)���a��F���:�������RX֪�$I�y����@���jB������YU�0q&��'%n,�&O�[�qm��YE}�:JUdX��*�|[z��k.�uk�0\�����"�x[���5�0tR#��CW�j�ʭ菊�	��t�'!pMdɭS3'}e�L����a�_~�v���O��ߠI�Y_.��z�i��������f�%���V���pw���:���Ҭ��u,Z�F�Ӹ�|��Y��!���60�L=Z{r(��ߒ�/��67��n=�x�V��4��e�+L��^���7�ݭ���A�o�F$�a�e�|�b�����28����m��>�榬�Qgǿ�Ԉ��Y Z�	�/��H�dE���dG��Չf>�Gc}�\	I�k[�?>�0�c^�R�?�0�%��
Mŝ��F���
;���Z�ɚIW	����]���S[UEw���[�:V{=�A|���f��:H���Ϸeav�XM'����|�3;$E��8j5�t���Q$����l���;-,Oz���(��ߏ+�7yR�_��r��(��=l�ϧ�:c�@ZA9���������b������骛���ֹJ���-�iV�e��k��gk�+�%�oht@��h�S������<�u:�n�q�[�u��߮7o�J���&��W�!�Xٙ��e/��
i�l�Lz��F�W7�y�������
�ឥY���	�_�[�*����5R\�p�f,I�b4�S�C��o��29�b�3�*죪�Ϩ��5n��T��P K]鋫�G/�S�]fb��䡿��gs`��ÏF�5Ė�<F�,�E��mN��� ˽� ��:������v`�]�_��� nR����ǿ ;6���?ΤčVٖ����e{�x\05�1gL�x*��Z�w4��c�m#�96D|hG�:fѲ�k8���mp��#j	D����ԛI�ߡ��EQ�ؘ�i�ո��=��Y���9�moI:�6dI*�ȁ�"O������(���'���Uq��7�/��#s�/�Ф�D�`[!g�肘�*�Ǽ�Y&n�,7�y7���Y��uhh�Ͻ��.������U+��=gF]c%5��|����䣦�ԁ�����x$K�[�6���cZ�Wώ�ל�<-)��|�٪a  +8h����`WD��ݿA��C��[��_�&ؒ�cx@�!���C��5b�/�@kX��Q�*��J}�ﵓ]��f�{���noq�U��;24����U�d��H�E<}���R]�]ޡ3��r]�%�4��^v�����X�Y������9���pr!����rB㫈C`@7�828Z%����y�1���]�2��ܙ��ӧ8��h�����	փOl�O��a��0�������I�g{�p���}	��V1���Cmƶ0�`�u��+�ž���]@MP���;�XO�\~���'�X�n�R����l����' i��^^�#�^�a�ZX"���	f# N��}��*!�X]}|t�"�z�*��f�N��1
]8�����FZ��/� ֨��`@t��A��������b|��HxL	n�S�Vd��e�%%%��t)B���en���/�F��=�4��'�f��A�#|Gw�i��(L|�~r֩}���N�5������槑�9�G�7�F���)>g��O��u[@I�k�7-���x��i�q��x����=�D]4mZE�����C�.�=���4L+�a���9
�6�P���W+�k���BEmDM���X�ؕpx�O��J{S+|LÎ��n���t)e����Yx��s�Rٲ��-���u���G�<T��Gއ�/��[�o�լҍ��1�u�o�2j�d��;�]?��t��k�H+�J'�z���B�0k��u�9��{Ew+3�b��3�m��I^O����@/;�ܶgl�!>�H�磔K��I�A^�(7��jQ�!;�&0���i�a�Z
m�nǅ�Zl��o`�Dg�f������p�z�U�"�O�k��%��Yg&[	b��٪a�����}T���ly'=��2�G�.��z�)�ߑ�1:+`|��tf��B؏m���ڣ#l'��&���l���A�,f"f���#�Uq�[�� \n��4�S�ssM>p��~BG�Py���Y�W~���\D���$����aQ�>�:L��(u.~.�N@������Tzr��<㋕�U{ʕ`ԧ�|?0��t~/��.Ռ:� 	��y�k��Z,��Z��w��D�0N��s)�=iB[.�S���J��1�V�sS�j��׊I��ϛ�!�[6��вz@�����&���7������� n[|���F�����6?��cG<_���Z'���6�(�^ǑD<�j�X�-|3
8����G�^\l"���w����_]���5]�Ȣ�!�c��|�$Jq�>%i��5��%7Eǝ15J��:i��$V= B�~���Hi��� l8��Yny&	w�e�΍'c�!�=�^&?B�"�mw�33�����i��s��g���%�2<�Wj�Z`u~���'�+D��-�q�4?��X��)�I���E-��i|�S%��+�r��`qs�P�vk} �J:�n��k�����[[�/��w�)�����9p�M�n��L�����2��WSl=	.~����&�(���>K[#�SO���]�q�<���L1	^rzg�"�țV|�Ӱ��#��'e�ʑ�?�K��u�a�ͤLҦ�8�7�����J���X�t��d0ʢT?�q�_$Ӊ��Kx�bRw��� ���&�N���G��tMW�<�5��U�;P��)F����b�*>&���il�cV2s���L;0��n�d%Qm�r������@�M��η,�4q��B�_~g�^\�	f��x�V���*�p�$���ʎ��Aq������/a�:�x׈gmEƔP���5�| Շs�̈Z$���zM	?�}y짧e�n���n�� ���HB��׹c^�]�*I�h5�.g[�Bwه��gu.��ivT����d<�0-�/�VuU ��C�?^����=?�'����'�[�����M�ͫ+������̒��{�nN�*A&��'������_�<s�l�}�K�M@A��o ���~�J��e�qB����^��=��y��M��ViB֝k�A���4��_���GS7�e円��<�>�>��{� !~1�H�`�_�(P�а9Υ�ٙ�9��t�J����n����B��è�o�TU��cu��Рgs���7]�QP�Q�訿�-���}g�����|�pSw�[W'�k-.�����I�瞦�.��G +�p�A�. �����}�oޛ �K�R�&���y<�����0kk��[/�D�*	-B@��0���>5�du���$�S~��/�*o��/5g�[�G��BhЭ�h�0�YJ?�tȲ����a�� ��U1qz0���D�$w�����<����.�]2Fy���_ZT�t�t�Au�Bg��oMS�q�������y��7���Zx��z�@��������νd�(�̼�pԢ�I�N�@��R���ɹّ���2�z�1w�2F�1z� �����	(M(���t�h=$�J�N�n�nad~�O����%h�����f7�B�ciQ�y}�adEr0��b��1]�؋�����D|�{[��$���*U6�rs��\#M�BA2C�c�o�\V:v�m�ў&IJJ�� zܔv`Z��j���;�y~��:H�S�ȍ8)=�n�5�q8&4�s��Y�?|w�+K�����ϝ*�V
���:�I�ѡa��F��'��%Z�"��,YY $Ȼ�'r�6�(�G��B���)�f�zv_Jό���w;�������F��%�ЗB�.-2���kNCQ��q
�_	'U���UA77O����8>TyOm�*���S֗��jA�P��-0��Z�F����QNH����\�ék��~��D��6��S��~ܳ�H�����0�p�,@��]$!y�O���R^��%�X3Et�X�l��XԞ��^9͞P*.��o����6o���<iR�4����o}�密2���1�B �-o��|үыjHb��A�T����c��]/�Y!��op�4��rE	k�I���\Ć�2S`���D5����$/��'����/�B�{M>����B����g�W$z�l
BD$8�1�:�Z�=��o���l�u�P��f��!9:�q���?_u���B-�mΛ��L|I�ܠo>��( �����4*���&TZ>�K��4�My�Īc��g�ʻ�xJ$~a������C������aBD�`כs��N���B��L2�y{VIT�,����t������eG�	JV#9
*�a�hG=�*��!�j�qs������-�!ۓ�wH�|wO�
5,Zd�6
&0~����ʅ�S
\��9_�?�&X������<w��uKM�6ۃ�=g��7j��ҝ�M$ 4V�4�F�D���[���Q�6t��'���\W�����;j����ѐ��wc�پP�׾O�8��MB#��J��f�j�j5dy�G��9˝f�س[��=��rݝ��HY�E�rt~��5�J���*1?G4_:*����������p���<��,�ou��Y��*\ �4!"vp�W��&��8#�V��(fm��l=%�~�PK��v����K��D�0{����ie�ת�<���eb����f �H��]��7e���g����GB��h����g�-Iƍ��[T�]�x�@[�R[�W����Sǻ�MoZ�&�7.�����N\�b�êUw�c=�rT��H��o��pKM�$!��ɲ�@��L/�ebv������-z�e� դ�!�J=�{qAq	X}4�Z��O���NDp�?���o�:bj~Ȑw�0��9[A<���fY��dY4�Ӕ#�zb��P�ypV�y�#a�̏��J��x��;����?k��I��R?/���ލ�POc��2T��=�&���9�)j<�1;�tj ��N�?���/�X�t?LR�y��7C_c������z�ʹp��L�ʌ�Ț������~�����C3ϺCe\ˁ`sn%u�xL�n�����Dx�fQ�};p��k��K�j������)1u��E[�����;��)��Zx����^�<�ѐ��E�kv+=S�q���d1�=a�ng�28�0�����	���8��>5���a�&�qL�.��7ޟpӵP(��3ӥ?+T<W�B��6)x9u��H�CK���°�u�6ܽ	��z�����+5�����>*[�ʾ��
���%��g1���y��s��%U�����<��Q�V��(�{~6wx��dόώ2��^[&s����C�Ky,��|p�����7?,Rˬ�g<m�gF��������n)�9h%�� q��_nU�66y���� �U�޻��е��93|��]>�A6O1͎�n�9e�Q��ez<އ��OE��3�kAXXT�o�2��9�~�OǸJ��W�{oy�N�KSML�!؉b=}��S���KE���џ��@�gȚR=n@�x�����]��{�{Κ��A,�>�&s��� ��O�7;�}��\����<��,��ȉ����D�j��9�x㣧��i����h\�����u"a��� �(��V��R�������1�.n�� @c�}?c���H����@ �������(�l>B��bPq��lg�툱+�8�����)K�R=�'9��K߅���wZ�B���T����J�>�xy71"��w11̂�7>�~$^_��j�BG4w��3��*RE�|ӈ�
���>�χH��b���^�Ւh��`��M�PQh���@�]ԗ��G�p5�p	�$y�D����sx75�P�(9!s�:P�|N%j;�@��|��,Dx�Ӏl��u~L�?�p�T�3Y���/V
��q����뾝X�Ϋ��exϸY�� �R'aQ�;;�Bl�&���g���6��,�۞�TSB���G�:wE=��i�����,�`ؐ�T,�#ۯ{�8���d����\>���ج�Up�b��>�ي��ؾ�)�38�w~V�GM,Q�=���S�.��um�Xvi_~�;`y�R����x@>�z---�!L����9��:@&W���r������O�i����t��Yg���E�AC���RNyN�.���Z�lY�][��aZE�!V��2$R2fJ���2�%��yC�
J����w]���sEP(	
Ձ�ɻb�J�a�q��zP���-Ň|��� ��;��Ѻ*�"�^���Fk���f� 
d��	�z9s�F(�\\\�"����PBv1(�=i���<�[['���h��X?!�`�a�<�nXn�?�+��gI�ob�ɲ�	Lg�Y6�����k��s�N7���6sc������+�v^n��!��"�������K�����F���	�����H.,$us�'���$��y-�$9��z/���t�u��e�K��,2�GZb�jn�_5���sRF�?X�ϟ����fR�;�*�L8�_Г>�w�\����ͩRx�pM��)��0h���]�<Y�B�N)0e>�� �sq�Cn&���b��9j�k�9���&,ӓŶu���#�?�Z�?)��P�+K�w�j�v����|�Y�Uk���:	��A4�]���2r(g� ���~�1;˩����)z�p�N̅�U4�=|��#�Ȍ�V��9)K.Ki�o�j��bS�����)��-���و��ʉk��lnŮ�[p.���)�T��ц:@���O��]@c��Y����������V�]*��-��8�)�Tio��K\�0���!�������}E��w��=�j"�W]�������?�<�y�(G�S})���9��6�&>Z\������&��J{=be\s����:Gs�X'{�F�^Nϥ���\�V�~=g<��w��}�����]��	F�Z�(Jם��"�c8)��w�Gq�.��۷fmEOWH\��5��<Dx��K���id�i�`v0ȐH~�����?��^k�fu?;�������5��;z�9��b��\����Ms�w��;N����Q���F���Z7�Nm1.�88m��E��ǭ�p� ��z\?N��csmqX��<���pԬG7�.
?��3�3�!/gý��F�)6<�B,����:�:�%���6��4;o~�q{۵|�����='�]e.�����[/B���F�����+�7�W����D��8z~��P�<"F�{r�E�L�^���?��,�"B[V��M���k{�Q|_v>�4�=Y
ן��K_2���G���⠹�����}�$�<�9NgrҜ>�|*[�8ⱗ���\����h��Y󉵰�BK{,�z
���\�����{X7�z�A��9G�-wU�)zF�֪����[���VG��n}�efu�Ё�;(��B��!r׹-���հ�\��s�+:!�,�*V��Z�N%����qxo
�hJ4�����z���L.���8]juGM��ŮL��Le�y;� O'J����~\�-�y҄�*kZ��XsXY�g���=��_dJ��i�E
�������<��6�r����r��T7xQPNFf�Ƕx��k�y|�~\>�{�%�}��9r���}t���V�413�;�Vvo/;��Ȉ|�	vV���Dma�	?�,�-pk��3)**�\�Wr�I�#U܋�{�Y0�GQ�K[[[?�>I�������j�Uk�m|�`��#ח�f ��q��]�ⶦ	��Z����t��_�IJ���#z����J�۶Y���� ���%w	0X[q��ȄSF��ԳW�"��x�'�
v���������{�w�4�x�t���Z+猴ܳF�}cw{r<�V�*3��`�h8����W��ӵh���sW�k�-��M=���Zv�+$�NR����j�rA�	Loc��
�Ə����(�;����D}���3k�Y�
kMp1�NY=llB^Sy�Ū4�en�E)���A��Ҩ�}�	q�kY���E��N]Lk�X�l$s�.<8::��(����=���K�C�������q��tT9M�"�*��1aĈ���G1/.|�cɩ&��kcm�[�X5�F���7p��+��\��t����7:oȟS�?T]n���'
(y����5�d4����ܖ��C�y���g�%��Gh� 6�2,k��۳����)��nذSF��K�x��,��H��\�� �.�l{�	��p���H�R�~n�����rlIRNG1h�7�sb�+��uH{���I��v� �de�`T���j�6n�����Ȥ��7_�܆4oA;Nw9���Wz܄��g�ٚK�Ӽ���y�Bu���e�$G�^4.�"��."b�%B��:������S�ݯIVs̽�iim�Ĝ��bBk�"[��O�1��o1�I�{�����aHwq��s|��-sG@�3�e����cL�����Q��05��u���N��.#P���3:{�����L<*����2zhХ߼N��!�F���\����x]����ɇ�|�A��Lm����cqB�V��bd�є�<$����$m�I���d?'����&���"j���`��1����OQ�K�`��\���%��M����s4���Ǥ���4Vc�ǵ--���r�+�Q�z��d���wA`�Ne@(�7ȑѡ���(۟%u������KZ'����Z~f��R��较B�x�s}�c�s�k�"wj7�J_Ǧ���.��/�kI��STId&|���9��u�J���f��\B�T���v�J�DAþ�yƤ��j� N&�ŝ�^j��NO��p�(w�{���tَ3^RCx!�������U��t� ���q�'�X �2p$���~��ӆhU�R��Ɛ*�O�efZ�t�W����i�4꨼=i��b��@k8�E"?���=<�*o$�N4��n{s��Q�mM���K����v�ræh����d3U��.�J�Y��A �aB�/�;�9t*�c��էMLW_���Z�@��n�95!*r��D]mm�|L:8�h��V�o�������-��~h���$�V�}���͌ڄ������ח!A%Y�1qH��"��rЫ��gl��S��Rp'���8FhI_ɍ����#���H����Y�׋���8�L0&��q��G�B���u�L�D���u(�������5~���7V*N{<���*I����8)J��4�r?ܶ�bL�IEY�W��woV�����]\Ȋf:E{8B���,8&D���݃�7�,��D����o�~����)u[.�)�c�M��4�K��"zB����:H�4YЋ4ϲ`N�����t����ͯݖ~*�z�<b��5�J��ɖ6��-��/RA��,��g��tw��d���o���S�L{e��������]��ZIp�<�&u�r[���Z��y�ڿϘ�
&�~��Q� ���.�۝2B�{�\��� ֖G��%u~��@�lrÞ���XI���×&qbP-��A��������V�(��[ac��p�+�"�ֱ$X�.�+>���)60�r�c����j�V�l{�Ԋ�$ ��<>�q�s#��:� �ͬ=�!����m�8���c�߬��_���?�t�#��j���~a����^��гB��;�i��v��?z�x#�ECM³syL���m%�C^��u��B�?���O>���Ů	W��0��n�E�wH��_f�t��
���.��>C�6���M^9dW�b�L�Ѭl��F���<N�܃�(�El�'bca?��a#	�"^5M�8ڥ�����8_�nv��E���!���7���l3����kK]�q���y Jje!��f�/���=����u�Y��"���#�F(ϲN��g�``�FX�"�A���|��孖��J�v���0�I��B��i���'}x�gX��E���h4ѡ�j�E���4o�O�rz��{�������@���r�3Q�)5Q m�ʊE�W�{3�V��[0Gq��0ԕ�a�R��̓
N����q';R�U�~g쫃C6f�GHG;��(�����Q�~W�.)�p����?_h�O~���E���`�3��ˎ���Q~1x��=~����$HLg#��zܞ��]�F�q������h����tꤨ"���^!2�7M�%1$�Y�Fʔ2š�����z��s��uB�}���6��qf�o�����:IDt��D�x��l��2_"���FV��*�����7�o��z�d�d_���j.�d���I$���"���?��J&�]����ڲ���uXGJ��j}��:&�ydV��6�QuM���Gx��BC�=l��(���-��hS��2���9�yD�̆�6I�͚�4���| ��P�ըOW�D�5��ߕ��OT	���Q�]�GW�悒�N�0�^hŽ���9����^�'!�������B�~oV[n���?g��*><��q~gE��ҥ�1{�WW�T�<�@+��ot�
�|��I2G[��Z���d�Li	G���c�:
'
3';���Z�$�>x�V�;�����| ����\h��lڞ�6D�9����R�����=ȎS77��e�jq2�Of��p��ޯ���;�d���o4}���K���G"�M�3.�{�a����=z�����F��}����8I������j�h�Ar䍻�����KS�Ompk���W��Ï��D6[�%ade���Q_���lZu1��E���]�l�����w��
��a1��؜C{k;�v���J}��Y��_ǡX�ѯw�$�����d�ū��B��g{��J|ۀ0���o�}QϜi3���Jo��a��!N��r�JD�DKR�|����V���Bq�D�Yֳ�jɚ'>����	iY��K�R0X����d��~|R�+��ڿO�%|��s���}ٚ=��y� �?��G�c�i������X�(M�p�e�f.{ؗ��(�ٰt��><_���]1,!0(����� �X��ٓA����?�Ur�=O������Wz5�nz�z.�@��v�5�]!�a	˗4��N�2��)JN��RO]TdO~�>\�A|�so�����4��Mq��,^��]8�>΢�f�����ǂ�$��s�E|�zm'�0�S�]4��g��7��@������l�K�ċt�'�v��ݶrd#��j.J��a�bv7���+��sr8��	u�����ڸ���1���y~@U����\6'ɏ�� ����Cw�s���0��5S�K�(yv�o�ML�}j)����e��+UAn�맫�ǜM�+[F��!;k������6*؟�`�p��B�L��*W��+�&��p�ϯ_�C�*����Tq��ClMt��-e�kϤS��1\T[fwgtu�c�GH�"�J�(:�C7���T��W${$�y���h���A(k�h�rB﮶f�A���矍Q�¨O%�a�1sa���`���c����?�um>��9\��;E��J��*�Ԅ�2� a٦��)R�'
k$v����e/��u��62r�"��P�:�Vs�	�FG$2QQ�Y�i�yr�BU$E:!��Q|f���:]|����s��f�����q���}�u|����,C������}zU�s	�\��9��m/J|*�����j��(6|���e�_�����Q��U�ϸ1O������_��Z�t�M����7��X"+�CR����s7�c,|�t�*�"�^���ǽ��X�K��l{�|8W���i�`��?6�rP6�u�c�6C-�?���7�.��υ!C��vm��	�B9sp�Z�b�q�'��� �����!�+�ytH;|l��*���һ�4)�N�w�ӱR'	����[���(ɛ�����z�K�O��?�@�`�t����'����>U�Sy]8{�ˍ�X@Y�]��ׇTmΰڊ�/�ܝE�y<s�Fv��c�=���)��- ^��9�b�e�� Y;��3�u�?u����|�(1s��<]t��Yg��_�i�O�]KV�,��"��7*d�5�?�o�Z�"C�{Mf�+�US��٧dh:��(ج����XA>����,�7���م�?TeN�I�G;_*!@\QKi,؇-7�l���w��ͦ��q�[H��u�P)��Y� �d�d�� �0�L�=�d�Ȟ��m�8�����r���~b���!!2���=������_�+!�g���oy�92~})����M��<�^F/�b.37������	������9�a����#Ł� m��Ϊ�(�E�8D\�S�U.��*����mۘ��т��N�$u�����ع3�y�P6@���)��om��ϫS�d���Hѕ�8�W��T����u��q�iw�U�QD�u-g������!�໷'&�����$t�g�~�r�l`S��w�f$�p
J3�F�g�녀�H�c�G������v^{���-n����rm`�������t��)s�쬎��xAL&��a�N���0>��̯������p���nVgK�t��%#D���Ƿ^_v����h�����/�J-�s���#�|r��X�{w����.��1��͟�h�W��z���e�d��M૸��]�uc�
�ɔ��Vp��u���֒���ЧJ�eɳ�h�������'���u;�0����Q�V���ΰ��	J�a[w������u��<ʱ�Sq�ʩ��(4"+����wg�DRl����U�`�;e���k�{���x�l�{�I���I'듨q;3_��7����鱒��4�(���j������!{=������%s`��KTug��-�{Rњ(�����p�=�����K�pX���j�qWA������&��Џ��Ct֫�~������h�<�s��9� �H�H.cnV��>.!� � {	7ec,Ó���al@�3'��R܉�;��������E,�b!"��X�ɛ���\-�o�j��Z������=<J���I] y����!YcG����9Ӳ_�ON�a [>V�X�L���+!��=�	�(U�:�p0�;CW�Ҫ��mz����V�n�(�7&����v���{Q����u�D�1�Cs���w��(O�C�c�^A�չ����?��;+7w�\�7oBE���\)�D��2%�s��n�5�A1�l��:
YZxA���c�Ղ<��7���ڊ�w��C�T�5����v^'�d�+l�]%O�sS��ս�P�ި90J����طB�N,�h�vɳ��K��L0�<�~u�>��y_@ό�5��$�����%���+4]�Ⱦ�݃R!��F���Ӿ�\�wD������6�����]�/�����17d�E� u������s����Ƀ���Ҽ�읍rJU�H"����1r+�ą(�8d���m������c$��͖+����D�¾��R�T�2����[�u݆+�LN�H�L��Jr�W�y�+���>&�gVZ}%?�>�z�\Dn`�N�2����!��A#��3���G����\�q�/��v�J�J�p������zȶ���u'�i�������Q��a�������j�z�u��}'�J]��l����[
YZr{m�+�]�h4r3U6ڱw2y�vny���	�Ő��X7֌p�<�����o�!{�r�tn��9X�`5���Qkv&)Y�����XA��: y?�A�o�,�,�3y7��1tE(�U\OM�E�[A�^
n,�����M�K�(>�P�Fz���Z�鋮y͏��5Lǘ�Z�8���T)7Y����O}%����F�60�_�3���V9��skS����g�m�D37f�-qmB��"ĆZ��_���.��"z����%랥Yi�.��^Ail�a����F}��իv���\;1v�e��L��o�!����Q��v��y��d筕�7�z?~y��&<|�{������Mw0��	$����M���Ȯj`_믁��FA�k�����3t�OA���e�(�w�;]y�Ӕ��c��{`692}���D]� J��,	 �DX˹3�f���9��N{f`�䌾>��-�������F�Ǒۻͧ)�{-±Q �����Z;+��rW����o�g�R��Nv���s� ��YK��A��w�*׫�����D?6��S�H��{��{�%d{+;��z9��m�t��U�jd��������-��K2'�����ٚ�p-]�nİ�����.C��㸯�6<�_=3�?O��Z���ע��ڕ*Œ�
=ht��r�-�m�w�p}�p��z-�p�CWeJ�j�B�����d`����ܓ��:qC]ݟ3[�����X�e4�o�oG^_ӓ�� ��s1-xݰӐ:pxprJ�� R�0�F��*%�q{�{�S�����uh}g�Zn��{g�O>6�hiߓ/��~�0\!�96c}i�������*�	�LW���t�?B�z��;q�Ĉ��~݀��\|4%�5���Y:�vԧ��s�Β�E���^��U�[ݐs,���>���v��@aY03@e��4U/�y��j��jb ��r&_�o�~v���|���*`�᪖�}��BV5�ǤK@�+��k�����58' � �9����d��pF8)�_�_'_�Zε��-�A����s�Ng��^b�O��Ԙ��^o__���lM�4\ː���M�D{��5��z��L�Z��^�����n]�O�{�}��`o�L$����5�`�W����E�H�G�?��z	e����|�(�h��	����(>cuG�HoQd?�A�����n�+���\C������������v��n���Y`�۟f���W�ep�'�RÒ�
j��>j�{b���f 
�U���N�Sb���Q<�T���@�k���F�QƧo�/�;��z�Q[P��j�&�>6ӽ	�A+��e]@O.N�h��` 
y����������p�� �ba6����%�ݔ��4��/E�ޚ�
�z��"���5���WjL2�˛ϊ��d5��\Dx��˂��a��1G�B{������T�H��j<��0�8D���4C��@�Ã�/���9�쥯��1����z�����q�%#�m���̜g\��:İʦVQӛ���w�*�%�	�Ś��ry yS�J��xD[J�^���Z����Kv��n���"�[=*�;��Sc�W����k9���~K��^�0k�O��ռ���1'��1�ҟ��Ő�J׬�l��k�ix�=:8�ŏ�_y|��&E�L,����(i]Ŝ�kߖ�䥩�ܶ�6s������;�� ���x�0��/������y��B�l����:�ɆQ=�Ō�f0w���,wm�"�r�)r�ss�KU%����!U�?�����_���zQR�L0�v�s{w�uڻ�%����������]D�jY��5m���Q�/�^�D�����(��>��S��ˠC��:V��]��e0m�,Y24R�#�㔉b��F�����h�G�yO
RD)����1�^��ॕ���k��.ׯm}���H����_�/"bQxm�JMIᗒ�nk�c���446q'L��1Ȓ��FΫ4�`��j1����+�S���Oa�L�M���P�Q���/���0�������R-U.!j���/E2����{�x�5%�`f3S܄��u��L���͛�<t��ggg�|���4V���]�t5T��!�k�A�νϝMv��u_)v��^���~>goP!܁JYu�(�)����[@=7�~�;f�s>��bv$��}��Ȕz�?�^�G|���#lT����X������1!b�U)D��ƛ݆�hE�0$�>�X�4Q\y�x�\���Y������ޜ0sC^(<(��˲~�n�FS��S��G+O�4;�{E�E���Y׃���"R�Y�ec����`��_�K�fu��Z�H�)R=�s�M������#����r��U�]3\sv�秳��z��إ
���-T�-���~��� 5L��[�o��/�����<�I�OGd���(�].xܺy?F��;��m�02�G��-�oaoA�Ӂ���w�ߍ�+#�n�����-"���]M��&|��!ZvhR�
[.^r'���N��Қ�����Qi� �^�������s��Wt}h9�Ӷ6�k�� <�#��3ٸh��������%�}5d LR�q���������r��o}*��W,\��:q�?�vK�$j�3v�9����"Q��_#�|a!��t��9��
�U{��_TT���,��~b�7���ˆ.;3����:h$�B�����tb>ӭv��vfS3��C2�P!�!���XqK��r:��7-Q[�/o9*�"w��ܝ3b'5R�����K�cm�5���9�_��:˄ֈӃu�3��u��~d&�rl|�`�b����Z��mKrwM�d��F,����mί�:�Z��-*�c������=O��ҟl��n5G&���k�O�i0ƕگo�R�����j]�fn��+�D�`��D��O�7��No�j�>�Mi���c��~���P�,{$�$G�Ǌ��lG�
��������Q�&78{�P�q��͝��{_���~���ǽ_���9^����K��k�r�R� 4F@�
�q�c6���e��j���`@�A��/�d Y�㈆�4x
�'_f�����+��ѷ��R���ܑԢr�Z-.���6ǻZ�w^j�+|�bjsg�I�� +"��٠1qgh~Y_$��w��=�lj>:#x�i�3����p�����
a=r����awF�!P�٢��Bi+��x�bd�z#`B�\t�X��U&?:m��djju�"�t�w��Uϭ� B������S�OvF���rNk+/oA,��o�7{�AU��v=F�)٘8>)��Wy�'"���W��eQ���6�堜&0��("����k�'�^=����m��^N�`�5��t.�ez�0}� �:�1�:��vM��q�`l?�z�3&���b
z27;�U�~�"t������wL7�	?c5��h�Ey�5���]�5�ps�q�[C�7�z-88�{@`��N��()��F,qᛰ_p�&�f��t����F?p�)۬�v^��%N�
.*���@=%���<��b[�C��w���(��[Q����ۃ{��8����5�nL}����ks��ppt[�U&�߇"BF�O:vUPg�	����m}
�=xx
��M߹���Y�0�{�]w�����'�@�xi%��^���3�>G��m[�\��6���������xT8cUd5"0)���OS�P��`OvΎ�����ي�56O��|x���9�Q��+bW��.�c�Z}����Ib���N۞��牄�y�U�RW�D���Ү�-�L��ɺ�67&	�
BwM��f�P�K#;�K#^T�.ff橄�׎yE���m붌���L�L�sH��;���Ҫ�G|�K��\���kB�M��j��/� �c%��͡���|�Z|�c�f�G�e)�<��p�������� ���[�%�r ��&��K|�tPI:�j9��}w�7���kH�{������ĕe���8AO��%}��x:�DRR�g��v��K�e��%4v-������(4>z\�#���r�bp���q���?�?2��cʭ;w�K�t���p>:F���ɪ)��4aq��G�D�/"JEg�F�5�`1O��u����2ɼh�\v���9_��
jw�,d\q�U�n��;� ˙)��CL��ΜivKл~����(�2x{,�<c�r�de�c����|��K?�M�f�S�l!����I�����х���_�U��N��~\)N0*e/#�}G���}���]�"Y�u��5�rR\�	l�u�ǡN�j?�5ߛę �`cs��U���xK���3�h���)/B&H��昂&A�NU�	��z�6��)��Y���X���JF��N�_*��Av%??���_1A�ߺkP�X�Y�]�*ZhR=����;�|S��EsƢ�8[���]�hp3�̯��f8S�Z'CW~��X`����fDF�����y��:?�#y�^�L�F�L�ɒ�~B���?�<����m�3Xkc�]6x�}v��' �:L�q�,�M7��^�*±�����)�mb�A��W
ȹ��0�(����Oޗ#��s�J������#Z�`z���A;�<6~�)F�*��ڜ�����$� �v���L/Ek�!e�Ҩ.{��ٷq_�B����	qa)|6�`ft�:iO�}�'%~>���� E����ű3�+���<����WY@��O�>��6.�Oz�7�H_��}��^��{�w[$����ڟ^�Vq�u��_�I�R�DF���kE��CQh|�����QL܃���(c>�B	s���+������ ^����܇Z��~�~4���S{`�E�(�#*t�Q��ʢ���^&�y���d#��El<
�i��xG�/�Z�0&b�_{�����U�1���h;�#&m{J-�Aޟ�,�M£�C��J.Z�1Ny
�8s��$5՞�@ϲ�]˅T������Ś�����(�V�ᜮOw������s`����|�n|~��7�`�8����cR���U����^j0_Z�TRZ��un����H�
���S��҆�k�)xa}H?OZ����f*��67 �ޙ.�B{y��x��r���:Ϗ>p`�!��:o�L��:����*QK�w�h�����[�_-q��U�!�HR�W� ��C�0޽�3���?�xN�4��.�����35�� 32�Ѝ��O�8�)�$NGV�\@�5����U������5�^�k����,��ٷ��~ʘ�5J[/��27&0��ǥ2��ON�+X��g=92B"¾s褂(�>^`�r��*Z���ǚ�|������$�ӨL�K%𶼾B���"�U�.�3�b4��tKw�Z�N�򭩈?������<�v�4���`���qm�Qz�\��z�����w�6kc����z;y���L�-���.��'KL�Ψ�8f��Y��Z�k��*6��������.����;��AmRW�3/58��O���q��$���V��&1q
$iM�W2�R0��V��1
���,>@��Z�s����g�/��E�·�*���=J(g?���#=b���)VJ����ˈ�z�nP��;��zqO�����U�������z����_(��1�٭�_�:O������?��t�3(�PB��.�?�@T�HD�&2c��R䂞R�*|~&�)��*h�\����߽�<�<"6T�����[}6M�E�`g����:`ܱg��9�ò�,�m7��ŔlP����u~7]$��L�<,����3!�BSZ���0r6�5�)�L7H�!:T��������gTA�P���CËY:�_
�Ҏ������x]�����,��)�/���WN~+~�+�$7�&�wvH$d)�̍�^�^��U�b]��&�p+����b��j]�v_S�,��=������"�K+����H�{<�l�ȳ��2�GS|ɫG�E��ڦ�k�nP���YlL����c%��޻TO�2����U �������J&�x�q���4;;c'���m�U?0�	�?A/m,���
'����
&æF�^��K���,���I��˅9|�#ٰm՗xȉ�=�J\�4�V�h���)�u�|�o��q�0��W��K���ޕ?Ыҷ�v�5�թj�u� c�b�6��^��_6��>�떨he�/Q��u��20:��.؟�[���o��qx�T���uP�#vǯt�Urs�B��X�n������<|��g��V���z���jp����/�� ��"� �͉_�Z�����H\���=U)#P����~Y��>��ű��n.m��i������c~aP�>T~�����"&D$C	hM�gS-	��%WG;��t�z����<K��*����y��������~4ӿ�W0���\B9��u�Wv�JDH���.n%�f)Bq�pw5�+��[�!��I�^�/�v$�o�ؒ��	�&ؤ�lT�C�8-��^�{`f�v��p�\��i4�d��z���\�d�����rt0�:/s�����!nY�G~���OJ��@ Y���{���L,>�b4+�������X�%b���>1�rD����%Te�ٽ������{
445模��/�C��L��R<��,*��)�%�u�%p�%�b�����:����A�I knOxnv+W�ݠ�<��;		r���v�ZdLV'i}n;�e���V����[$�F��Jˎ�l�q��e�LH`E����b���W,�x'L��[Ak�xy:����Z��n�⋾��Wz��f*�!�f)��t�c�����ܫ*9ε�]gˤf25ă�c��h/mK�{<�{��'��9�Z��:�9�:^{�솿0�$'MCIi���G��|&�8s���b>����l�޿�4�*#XJ��0���\uF#��=�[.�ӼW����ٜ�_y���c!0	��:��&��C�f����4�_:�����R�Q�!/0|&~��j�^ �K\z(��Ԓ���E)9E�?~3���*QK�P�E�.�3�/�2��`8��-�#9E�Kz~�g�� iIڮ�f��-��Wb
�uS�vj�
�XkO�X'ݻ����?�#��	 ���2=NN>c�Ab���~�_i,qbRe�e"J;V��d�J���e�.�o���ުI��7S�c�h443)��r++�u��&�p�ґf�5fJ-
w��KCo�AA2���0���t,y�z��t~Mn�\��ӽ���g�E��LGW@��e��۴�	CM�Z4�����&��~i��.��4�3֦�����86�X,�=9/zC	�^��<���2U�O���i�Ğ �����IX�^��]������l���M�E�~�h����G�ZP�T�׬����L(X*H��mQr5w��J�P���\H4�7����1N����L4�\���k�F�0����:�s�W��,��k�?�f��J7�П�Td���D�0�'��^A��2����w?���n�t1x%�VѶ`V���~�ʕ�{،�TTUZ�ku��g����E_�2�Ӹ{�C*�+I}����J#��ϑ����ɇD�*a�wp�>��q;=+�6��PSU� �{��L��M�a��'6�[y�T)�.�}�%N����)��(���A�4���[zf|���໘�A��7M�$��*��:8���y�*�%���uXu�WOȻ81�%'C#�Z�m��u�����~�]�p��
.J�S,⳵�U҅<Cb2Q��������bn٣��Ɵ��:6�9i�3e�S'�CDYbM��S9S�����1���I��وG�&[�V+�B�?�����A��pgB�v�>�Gƴ�Q�BnΚ0p����E�2��I������X �1m������adG��	��i�!��~�f\Ԭ��w����g}	?~z��]�8r^q5"��S������H���+�}�)�K�g�ӯG��M�W�Y�
�L�~p�}�j�;�U���(�7�\�C`�->˾��w���ƻ�`��o�E�i[t��D���P��Q[�7ӭ�$R�T-�g"PDm��$0�Ǐ}�R|z��W,�'ф��%=�$�rZ���6�B�d�G�ezQ��n�҇�>ɚ1נ���A����x����&�3�1�ͮ�y�%���n��u�Fw͔�rt�3[GRɄ��Y?�@����ٓ0�}\�d&��j�S6:0y��/�]��6����l�;�E<DוM��s,�O��(3���v��<O�����<`��<��mv�\���f�D���,�2�]>������<'��>�gee�x?���8�D[�
�9	;ji �c�<t�B����lUJƚ�R�/����jg���͈MT�!<;g���/@�A�Ģ���<CKɕ�gz8�T�f��IP�}Mbؿa�s���|I%4��Ϧw��Կ-/ȳpGݷ�������s��x�3Kk>�LZ�Ҽ�x�r�@��^���t]J��{v���P������L�P���xX}L�VQ�c'���`�}������3�a��O�����o��'�ՑRJ~í�@L��`�!�(5�B����d(װ��%�H�Zs�ʩS�i�(zL�̲F8�6�$��^�3������LNP{�6)�\�X��P�wF����ȁ���|��d�`��H��2��7��@H����|��8nHПB�|�k���A��� �nl����o�X+�q�*��-lvy)�GJ-�
�l,�r�6�[���S���ZS�z��^!7ЪlO_�ӈ)t��A��/ʞ����_��|$�;j_�F���Րj!��k،CH�H�c�+�r���i�T��P�嫻�c}���
�>iY���Q.t�7�u|��b���#-cp�kTϠn�,������Ծ���I
@�<h����}��go�D�a���kk�d��w6����q�����6�U�+o�FWG�a�]��ۛ��b��0��[2���>	�[�T� Ŀ��?�D�k�YzMV����v�9M�����Bt�𲊊�o�y.l��9g��V��Bg����n�K�%����ӣKŽ"�#>od�����X&o��[�Ք�T�&4��X�8#����/�F\�Hiw��_Hv�>]���������dm��;:B��.����A(eE�_�Z�2���P��xQ���v9W�]Ffk�
�1ͅ3T���(R�O�]#}��n���)�k�-�w��YC\"AK����<_��m��T���xBʥ�ndH���O~d��8qt�Q7����n���[��w�u���X���e�l��zJC�W��V�de��[�=n&$�����msF�O�[-�8]'�碔:�j杍b�g/f��"�4�t�kBc&|0�Z�#NS\���3ӶN�!*�/�9%�ۅ��յ������U��u����Q�e��	����,+r�h%�Z|�L
����e��Z��_ؠ�JT�Ko}wI��7W���		�W��X�Qq��~��Bnd"���s+5�~�0AK�SO���e�!�Bc�'�����Q�#�F"�n�lo�U:Ϙ������H���?�y��q����t!lS�9
q�\N2�?�_YW��$������Z8�����[����^�A�!��~(�f�ؤ$�Ms�2�b�p5�-M�O���-h�Sud��9�-�HX�����+�f�ip���;����;���'Hz2l��ى�K�nݜ�!�3:fO-Fc W�DbZ߷��!�W�m�.{
�ʮMQ.gr����߸������G�;>�(�H��KMO�/����:w�Zg�W�����d��,`����;�ԏ-޽�?p���`�Ǽ�wGGd�c=�?G�G[���������\s��>N��sM�
�U��7S2Q�~hL����w-Ż|�'�^(�n��͢>���VnU�r�H�_0����Z���s�z��Y���HF��'��f�*!Pj��戹Q���B�<������:=��A���Mۘ��������1��Q�p�(W�d�?0)�N}Y7��3ڻh_�,�]1�w/�S�O�1�y+:񼴊�9�ش��.@�m��\*e]����m���.i��@T�}o�DUF莖Y6���vp�H�����B�f�kQ6p4K��ZD,ېm���&,g�<��}�FG���I�O�����[���;����<#t�c\����S�t��hm�:ky��^0W���H�$�ΣΎ�����@�*�������I9J��8,�V���Y(#�_��#�P��~�Qw�Wֽ�-�:�cYgh��h��Hpl���\L^y��B����n��>Ș��$��'��7�8�j't�A���zA�x^$����g6�@����i�e�I�^���q��]��ǫ:c����UI+jQ���m�t���B8�����R������z&y�Z�0�Cjd�V{g�?=��.�q�TkSX���~I�":��]�����4���lUn�v�����~��B�g�̕��5�57�Z�fF7���VTk�3�,tqK��ܸc�}��xS��>��n�}>��H{3�����J���k��Oh��]}��D�d�ݎ�<=D^����D��,�I����<9�<وQ�>U�j�\6n�I��[4����`j�t�O7�ձr�|��j������P�M���ۻ��7���I,��ׯwI��|����2�܎ưX�Kم�o55/��&�� P_�~tTқ�jl�^f_�>�>���ע����S��4~�p�uM�{�+MKP��z��0�>6����^ŷ��{O�&���ϮlQ[�ڹ��ͺ��h���{���%X����^Z�ܨ��SEc�Y����q�Vj���ՌC��/,1e�dD�˙[+U+ˌ�A�����3X���_�ZҤX7��CZo�nD>ŭNp4=��/��UE�� +o��5vr�ן��3�O|irE�nmgNj�.n�z��@��x��S�C������X��)VcΣ��k�mn�jЀi�R�]�T��+&|��h�d��������\u�B<���;�vǬ�LS�K����OhR��~%�u�����'��)���L�����OLd�Ĝ|�_\WB%(��О���.�殛'On�1�>d/~U���:�}��y���	��z���(+֔M7Kǀ���/=W{v)|f���l�&��!���g�Q�q��ɵ��w�5��h���2�0�qb�h�V;��[v���^�w�v�KS��3���	���60��=�$�O���I�w��b<�}�,k��S�L� yUv����#��� ��a/�wV�M��2�`cG:X+�_�������PF����v-��p��Ȼ�N�$N`�n��Q8�;�A������=��\������}�MCC���F��_L▨��β���E� ���!����㎎�Bk$�5��`_�kaaa����@J��ɫ�������`aU?�Z��/���IR�l�k������P��p��{�n���[Ωa������u?�\��G�Jbe���M�z(��*�˖���5��LqeB<�,��/+��٧����	�������L���8$������o��Oq,I�vFu�LB��<�ݲ�@�_e�I��a�U͑���wզ�{��S#��;�캎���>k��o�F������w}�(�>���11μ�8{���
{�e]F��7�ag��X�"ʋ��s?
����_cyn}/����N ��g�Iq�����/����5�^Bl��ޛ׭�b>�ǟ�p�p���U���dMLpQ��JA�=���C�2���U��9�>�$�ײ�ob @g�R6�n�w��,���Խu��v�:�����=#(����7��|e���
�o=���:��I���1�G�#]4cS�y���̀:����+��ѶV��*�rn��i�%�^�[ �AEW��	V��:&^]N�1���l��Xκ�FO��>�V�~�ա77K�Q�,��7���րs���G�����*����1��v��U}s�H����	u��S������RiG��j���$X��LÙ�wD9�s$�?�T�xSj�޺�	K��~�7vav�����~b#��nŌ�u��������K�!���6�׺V#9�o��e��0c�>���']�u���\{l���������B}Y�k�AS��B��F3�ޖ�\)��Ҏ݋[��i��Y�5��=-�G���'Gʯ�9�s�eB�c�FK�K?x��I[N9Z�o7T�d[y���͵*��]9h<�K!���	�?�fF~E�Tp��s�ظ��X���;U\��Sv�7�7��ه���;z(p�KSn�����<�/W�m!w�y?��J�ȼ��v�����<��0�=��������dGњBCㅫ�%=&���:<}R��$N����l0RQv��眿ˏ�^i]��R��t��^�4�]��3	�K��u��)��ąg��y����Q���X	ON�'�w�"�g�:��FWVƐ[����Xb�yQ��ҩ���j�KV��D�ڌ�΅ɭɆڙ�W��6�pZK.��ry�p[�[��*�eLT�n��np��*������µ^���?N��岒�!���%[
�����\�{yC�?��R����L���]��O�U%�Y����g6�.")�aU���m�^��K��F$�����p���������Mc"<O�ɸ��:{�9�*{��w�b�x��<�)╩�����!���(Og�<���aE��]�0JS����%oF�`��o8(Z|u��#ా��6�R�8�LMM��Y���[�mlX����['UoE�5\��=2�e3e���:1v��c�3:�����ks1IC̠�*�8�ޘP2�g�kФ���M�Ԑ��v�t�tRu8��Nlm�n������F����΢��N4#���B͵��~�!:�����f:h�2Qw��|�'������i9;�h[CI�����q��ӈl��}����M�z���H��*��u����H��brn���;�~�����+�̋(���<��4��Dy�qǎd�
��-�u�z;���'_����i%@I��p����T.E�Y_����#/|�G��+ꎫ�.zډ�N��-�-��'�#N�ǆ����}IWt᣸���*������[3ʃfd���«��iae��
t 9�|�	<���ã[��,<���.�.�5����7;�N�]"����<�N�?��V%:^�U��1a܇>�k�� cBr��3jnH����E(��]<�[�°.�J�o�Nxa�r�V�ت򆠡��߰��u��
x��[=�D�'��GGzt� ��>{���<���O8�-Ğٷ��Ϊ�yK�h�Cj��X��7;/n���(��x;L���  ).�kŬ��%[V7��͢q�@�Ѯ�R.�A���kllM��$>N֗�a�G�'��'�����������Rc�Q��)�; \[�l������zK�4�%>t�l]}U���l����5��b�=���H�t�E qg�Ýu��hc��6>ԏ>JD��o�X����8ʨ4�����[�*�D��\����\�B|ڿ+���)Gue���_��Ǘ��9���(g��d��#QW0E�@�{p���m����.e_�?�Ԯ�<̾׎	>*�c��aqy}��$vi���1
��0���V�ޝ�C��ЙO��s��]���LqIm�dۆ�UD�Tu�po�_��dF݄CY���%��{����������ki����Ķܛ�8���m��{V�3b�u�r�N�������zM��dz��$�͠��%JZ򺤅S�� \�m46lK�]���A���&�%��_\���e#�D�n���F���m�~��P�M�)�b1��������&J_���Dr�->oo1�<#.b�q� ���f�E��b�0e�8�\����;�Q*��%O�v�����aS�"o0D� j$s�/�}}B�����Y�	���_�ћ�Ï������}�D�PȐ�i�m�T}����&%4O�!B@�/�{�%�3�D�����
!��� ��0�xf�����	���J8�<�|����NA�+�ؚ��g����Ͻ�����:6�׀�mu�m�j�#�T���;_9�x�����P�-�jh�!����뒻�X�A����I#CY���]�%�B��1UJ4\Z�c���Ո8��"�$��sgy�_h�4��U�&��ϊ��|�P+�����͇\�F<�ے�?��EN�sQJu�t"d��d`�qsrОk������.}�.&�;�&�(*v;_����n�Ϡ��%!7���*3���F$�	ߏ]���29��?��B7��՟}۵�W>���������:�)��eYdy�'�G��Z�Q·������w���ƴZ])
�oݵ�Q�z�6t��oߘbۑ������O�ֿ$��l�-8�{_eo���vx|�(kM	��'�]�\0�ǍjL$%���]��T�cQ6NF����\+�w�-g�x�_r��`�fG��l��߆n�'dU&�a��ٽZciI�J���Jۂ�Ș>�]�C���t)^��sjs/��"M$�5�(Ux/ɱq\S+XELMP�n�|9m.�\����-�f�+ rw)7�z�;[Dd$tu�T�6�/��Wڇ�(��i0(X��|����/b�a�g�Ӥ�^����U�G���L:z��ç^�>���3k0����
�� ���%��F����!
M�?FЏ���+�/ɫE�ql�<��4�o� :�2n�W��H$\xX>T{���˼ǿ{`�>40����\�fD����HL��<��=�sz(���MK!�s���vaycK�f�.�据�S��
�{����hm��Hܺt��]Ϥɿa��@�(���Ӆf�Z���ǭ2n
j~�;#q�$���D�}<�{g]�"j�r?K�`�x�~8���"�\����
��bL������w�������x�L^l`����nc7��|/����>�\�܌�K/t�W���W2�x����ݬ2%P����1��&�P��˷-�cy���ê��&a��"�lO�Ѯr�m�Ye�-�HTR;̝����0�k��eC�|��҈�q��<��P��p�������a)����=�����\��5gW;��I�x��oPo{�|�U:?��I��=0��}�ECp�b��u�bɀ3�&Y���;��z�������xN���O����OpD<���P�|�9�I3+��4b���j�[��%�8#R��%�  C�,Qn*~�AvMM�RRU���^^2�u�9񎆄�	q��/j�#��EQ�o��:��SA~[��1�Tt\Z8�i�J�Ã�+jjs��Y{��c�W0�r�Z����oN�e�������h��k���/>>K��f!5*��k�`�PI������Ơ���u��C7=]o�O�C�l �B���^���lr�I%N��W,.k��kPRg�
����^O��㝈�3>X���q^�B�Ux�͘����U�>
�����h�k�z�k�Œ���S{q/�,�����a������:�1�AH�b�S���-��W�erNghNWn~ј����;�X�.;�r֐,gIr���O�Z+#`��!Vn�8م�fg2���������%e%���|oƋ;/��R&�X,�=E���r������$��<���s��{�'h�2g}<�����6 $��Oj>���:�������׆[��1�~�� �$��,ʪ���[���<���ݚR��:9�����m�'��r�8Y�HJ�ƾ�\n�q\�8�#k�Qh�֍D�.�BN�rX=E�$~��-]{�L:à8J���Nk�Ew�ID�%�0v��g��;�����J�lw!�M��#��� :�s���E�;�g�mW�5��뭜�|��kG��+s)H�+���<��:����*��p׋ڤ���h���%9�:?6A�Y�|!v��}��v��^=�����7��:@9h�Z#_��<%��Qg%��(�ԭ�*j�sP��o���o.��'8��'̷ߘ��0��e������-����V5���> *166��ge}�#,,�́���<y�9��z>�IȚ�m�9F  �J>_�M�TC�3�+��a�;[H�s@���7��e��T�r�P����/�����rU"�h^� ƭB�ؽ��簀����S�ɝ>w6�0���:�K*\o�e���>����2�	%�G0��ҍ�?t���Q&�N}����1L��Ŧ����T���ᆚ�L>����^?���2��_j��i�߫N>���/�N�x�uv�V�NA�g+��{]��� ����u7��3���t���I��&L���.��������`��/m-�a�%=�큡�8o�뵻�a���㑬�@י��&iiIh�^X���OVso44�%��M��2F^ |zrlp��"=���pJ
v[��N�t�0j��M��f�0����� �W�Ltv[�!���).�ɚ�n�	۴*��[�+"��v�1SI�L��ص�ʯ��&8-�S$���7_�6�t��Ӏ���Wy5^��\�2���*v7�/���?�h8��������byw���I�΂��v�	ֶ|̈́j���MYgb{u����U�~!%)��Y��t�y���� ��5�Ny�'݃qq���z�5P�4�4=�5	 SBئ��/��aEWF�_��i߂2tm���:7�sff�]�,|�����-cšt	X8~�����Cw?���QF8U����L��J��$����O:�-��e��4疤��У(�J���1�df��	�v0N}�,�VWp�|�ݢoi�@�iQ�8]F$��S�b���<����]�����dU)����1|�1ǤJdd�I��aУ�����M"��C��L�V��{�e�D����ƶ�Ł?�D�u# �#�w���Hۦ�û/��$��Ia�h��6}qN���+i���A���� ;=mqQC��+��~�Q.�S:��W���­n���%�1םlp�����C������q���" �齖81���/�(��Ay� �}��w�G�!QQK3��f�bͩo#��;��n�W�5na�<��l�>�{aռ^��8܌�'nXO����cN�/��w� י�h�)hc����$��Q�i�G.�1G�j����KS�]ryE���ۋ��m{h������+Jd���h���C�i}�G�ZR\��+�ܙ�+���r�9���r#0YC!&]��W˰?�K�]L8V#h4Cjˎ78��N���3�7�F��7�&M`�D�3x�&K5����O\�B|ef�|��qS{�5ccIeݙ;o�gbV�o��bŜ�3�!տ٩u�	��P'��y�ߪ���XO��;����
�<���Ӱ@��l��}����ON蠒Y9!"����4���r}���B��{%�<�Dֹ	q�����5�l����m��i�?}b�=u���ϡ16f[�艔7���1ۙ�ƙ�޺3�n�71}c��ڙp��* d3�{A�]N�w$�t��!~���=H�t@ۨx�����`Wr���{��z��8��8]����?����ȷ1s�
��V�VFk�[0<T�0I��*g�z+r2 ��I����%��4#�8N��\R�����K�Z��/D!�;f�$M�\P!!a�ЄT>�Ȃ���{Zg������z�m��ڌOO��-ʓ��*Ch�����=�[��Z�HN�'0�d1?k���F��;ߍ�ݕ�bv��SPF:�af���oYZ!@ȊJ�Y%Fά�v� ͤ�n����x���_< �kĵ�\���/�9V�Ky��o�z�����wOS������o��3�Vi�������'��������G c֬�+�sqW�к�D5��n�e݇��o9�7���\9:�������$���<�Nh��o���C�^���� o�x�݌r�Y���ַ�g��K;���s�,&i��i��L�D��=3�w�F;�ϔ]O[���>�!<f\/��'ػ���o͑tA�-��h�6��x�/[>�wvA}���ge�p'K$T)�C�,>oJY�K#a8g���h���e:o����]�����Ŕ��JT���8����H: �ڞV~ϛ�;p���n x���&G�����������"1}���Nv��Q�����kyt�4S��<c']���5nn�;�W/[df�����3��R��^���+��� �0�	(��E,qR��ٝ�pz�Ү�
pX;l��&�(s SG��� &�=�;��P�9�7�+�8���ªV_�VP0�2}ǙR��8����H����[E\*�l�l���_n�פ�A7%���㫞����g_}�]��1~�����	�� ��}�Xb!�&����NDo�����7��X����;�~��A����"^�mk��e�?�X�碌����98�By�?�b�g��1��s��v�6��a��-^rh ��>!�RF�"@�Tj\���. 6.ކ��S��a���i�@��DV���~��g/��n$��<P��y�q����}p�J�K��u�AE���VX(��"΂~1��1�yf�>HDAx���l�$Df�,*�%*Jk"��e2G���3�	5���1�����*��e�x�=�׻hD�74�ԇ�<�C��2�B�ԋ�@�]�M볁�4�In;q���t[w2 4@�(eF���>=@9^�,_�{��M߃�O���y�Ω2�C��W�s���5��~��
ķ>]�I!��	��a��D��V�t�R]%�Wh�`�'�AkD�l�#c⹻e�\NS��2�+Q�M�
wL�lB�γJX��Һ�[�)�@��R�Z�>�L]�U\F�fF(_��D�m��5�s�:u�qq�)l�5�9AR��#o�A�����tϸ������0�Ah���<̡��T�$B����/�%�煡��������'[ܰL	����	\Jy	��n+Q\�?��g]ol��[�Y)J�\�hF��d���	�g�mD'�G�{xٝ���vN��_J2�����\|0ש��ԓ�w�`ΐ��㞧�%�1�|�jm����@�_Ƹ �[��C$E{�=�57^//�R|6r�a2�ϋ+-
� ��F��	-���i����P�b;/��W��6��㹔#���:Ƀp9 ͒����0Fmf�ώ"􆈐1�̡�[n���e�5Q%��
��9�=x�e�.���IA��Ǳ܆uwK膣Ezd��a�w�l�={��YӍ��>L2�z�xl�|D��i����%,��kv�QG��t���n��J)����`��l�n8e�Ϻk�'|��ځG��|G^[Ա���L���އ��x���m4��(r�xU$��O��A���8'�ثD����k��?@҂Y_h<�!4�Ɨ]�/V�+g���>�4J���J�}�x�VPF8c���±zA��̋M��g�|d��d����~FiL��cA�j��%�@>c:�+��Fk�0{�,.�ֶi^� �(y����>p�sSx�=;;���yѿ3[+X�qo�Hql^�[o�gvGN�uM�/��f}���Is��F�*-S˟F�}�H�k{�}a��`"�d��OT����3��A�hy	O�;g��ZlS@�D��Q���;%bo�6ƞ��hg#E�U_��F�A�tH7�)
H)�).H��(]��t�t#���� -Ͳ�t.������;�2���>���|��y^N�:>�?�+�mi�|��eA>TߠT��~0??�̟�o�~�	��~�>�������d�;]���W=���w����Vɳ�zKs�_�F�,~"`S��u�kRA����4�5>���%	��_���~b9�+0_u4�:8�h!w\������c�졏��'�e]L?K\��5���vN[<�u��H���ʍ���{�gU�L���b�PD�#V�	�9j1�F�|���qv̛���u˪��Of��fQ-Q3�)����QJ�T�5�t�lR�]D�`qÝ_�Vۗ�O���,n��X4���u���	h���O&	:e����JZ�$al�}g�H�#iQ��@��3I�����F���&�7�lFq�	g�5j�Ky��1�&�z"����
Oz��^(x8�%� ����+�M���%lm�}��N��w�ҍtw����r�C�/�q��̖��Gs���`G�k�u�!)�V�z4�����j�%��+�д��f��/���j��K��w�����nj�l���ߴ�����+�W�x���2/�p�r|�=a�b��'��g�����*������d����o*�d���x����f�ec�
`0F@���]�_cZ�i����=<���$�	��>l+}����7}�u�퓍�U��(�.�OO؞����0ER/�`�0^G��,���Oz=!o�X1��r�z�g	��ڊ\�����*k��K/K���/�g8�����{�./O��O��`n�&M�ۃ�+W��ʬI����B�0� n��+�
ד�F���ʌ	*�~��3O�/�G�J	�1X�-�����A��nͼc�zXF�i�7�C2�/e�6���N���#�6ǸfS&�_9K2*���9��PU� ����pA	��oO��
�6wB7��xK���3�TjĊ#��0y�H#*�[����.�V��v]�x�>r�Ű�w,L%���G������*wh�QĜ��i`vl�ߛg�k$�=	o{�֝��eo&=�.�g&�Ұ�l�lﷵ(/���4��+O�0l�Rݥ��`��$S�V�<�LtҁtWJ!�f�9�o�������bf�u�&��kjK뉢�̡L/Z���0;��L��������+שmwZ�2���4xl�;)�8{e�'j ��ۣ�M���:=�.T�Ѐ��H��0�.��������1ܗ�L��ó�?�/�F;׍��J�iᗕ͠�M�
��-��J��	 � ��1J����ܢ��NJ%Ծ��4M��`!�>�>⨞u~қ�)��S���V@tt����:��'%%7촋F׷�F���}Q~@W��٠�lXǏ�A�Ȝ��j.�Q�'��y�����'%%a`t)���	RNz�1���?n�>��*v��b>��� �/��1������K���l���p}���r�MҪ��؛�-{�9�R��S��﬎��Xzׯ_�5]rH$r\��֜Q���v"--��2�Z���}P+n�&�=�U�bV�}ʫ��yN�7��zh3�O
�Z.�:��̗�Gmٔ=�D��o\c����3�4���18��;����o��?�`��>�>���B�s�(�]����ǃHܦN]$��R���	�!Ѓ�RD�G�/q5k��z�$�L��zj�3�5�t�%**ՠ�}�ֱ��8"˞�c�Joo���`8]r�E�� �v�e,t3B�sn���\Џfu��ҨX��9�0��>=q�Oc��7��/�(��j?r�������I`� 3L
��Sϱzܵ�>n�
 ���'ω~h�9K����$��yм���U�e^s	����,�b��u�+�G�Rn�<A�m+�F�V�3R2�9D�:��̇�������桁�\�G=#��R^jglKn���w`խ���+����w�^[y|�(�SU����������6�����+���er����7�.�&�m4�wu�5M�^� v�I�((��}�ޣ\���=n�)���-�L#�h�dۋG?\����4�4O������
�	�*s|Q����9��J��~:��^��ߟ�Z���$G�G��]��Z�.3�E�_`����O���,�PN$=��,��4P��y��u�K�~�;(�|m2��|!qT�!_	�gy{7�� �^:�1{`�J7!:��'��\T�zA��İ�����/�N��*�j!�&��xG栗RP��=�=#�aΣ�W	J�۫NT���Y�z���hr'/It�J���T�{����u��@j|�;��N��b��S��?�ң�?8��f0g��t���%�d�s�$*����ћU���B���٭��?����5���uӼ��ʀ��r���W�Ύ#9&��ݗ��]�ß(Te���^���qG�E`T�Ys�Ik�Pgp���B�L�rt`z�g�h༖������ך����3Skf�ד+�g�M:rHZ���l��'sxyw�5��< �d�&br��/���x�߈S��Ⱥ��Q�g����JK��CV�V��)��e�u*�҅�02�a�[0����c�n��hz�|(��@�9�/��^X0=��%���x������.a����m��UQ��&0��?�[�yy��� ����	fMϵ�ټ��<ݩ����]8�Z����������fD#���I؁�ɺ���8+nӆ7�X����α z����D��yL����L���ͪ��S���� ��������(2NAQ��#_,���Z1=e%��;�QPS�ۯo�@֤^���Sֆ�&l�(�+�O����hf�W1t�J�������SW��-�]����_4Н�a������"��/�;;Y�C��4��0CTf�-���-%��L����ϊ�`�.���I���G򀿖N�>V��gK&����4mx�x�j���.��5p�J�^�)帯�A�1Pm�?�	��QjP�֫���ο1�4x���|�?�d��&�V��cA�M�IR������)����f��ͫWM.	/)�<znӭH�uuuj��[x�����OA�WC���˽_ ���lf�bIX<�_~��
��������t�)�b�T7��ñG>�{~s7}�1��b����W(�+˿["8Iq��h���	j����n�����@M�/��c��9�*"}�/��jS~P�8�{���r��o��
�K��^���ٞv�K�Z�׎���(�����	$�ڟ��6�_$������	8��TZ�d��z,6Y蘿��	�#������kX�BЗ@��g����=_�0˩�p�KJB"y�/����D| �f���u�sj���t��s)�7��U(:�֪֡f��ww���M��l��?���U�>��R=�~x�zG��W��~�d�e�ե���s���6���y��p���d\=QB�_B�d#�L��3��]2m&�i;~��2Iqѭ˴�D$$p�����i�&UC3���.6��Z�!�હ���+�v~�X��o���O�N �P��K����$��&S�ne��25/�v�$�q��az��ʾ�d8eU /�iT<��bmt�%H�M�����Ә�p%oP���k�|�8���m����qS�4H��^��bLb�2��Tط�nX����?�u���z\�Pe��U�<�Ү}��DZ���C?v�*!��4̢t~j���E��O�?���2tG�F?f�T�avW&��\%��B6q_W�L_���B�ޢ���ۈo�vj��X���2
�u�x��g��ҵ�ǷL�C�sS������q����8��|	.�mX���}�D�u��Y���mʃ�K��[2�d��>���;z�J�����?7;�%�htf��y�j%����=Ce����E�0ڳ�clek|��J��b#�m��ҹ�����A��]��C�[��sD7��j��;�)H��^oMb�����Z��w�U�x��Ȅ�fP@`1;�L}��mp7�A�����:Qx�9~��i�8tvLH�˔���t�P�� ��)���Y�㍝�S��ț�N"Moӛw���ulm�"��>k�x��AgOlpr����I�;��u}�w!\*c���.�(~SV)1�����������t�O�V�a���`��8�����,9�+����z����sA"}K�n<pd}?���Rz��!�&�t���b������So�ĢP~���ë>$c��M[�R����=���k��'���G�`�bg�����\i����B���Dڂyn�R��2K�Ϗ��Vwn�����2b�a+�`uˮ�o�$H��������ӾR�ܱ�D���$��%��G<�R�fj-���X�-�RJm�H��{��8��XI�$qj)9�A�/�~+�(y\2Be��=��@�5O��J���/�9$wq`�{�-����^���0�vzv6�{{��+�I�[�rE	�y�s�Z�G7�z�$�[CXgwQ)��C�b���B�����P�u�%Fq�Ge����)��usV|�eCRB-n
Ov�ަ#���y'O�}��	]v����%a;CD>�S��[��3�RN�!	$�:����XR5�\vI\�t�/��*��A]��<��}��Ŭݞe@���_Cg��l����]m���Z��YA2�9:hZ�$g��R�47��5��(.�@�XtJ
~��m.���s龺ݹ��$5���\J�1�Ҽ#`����n�K�V�Mq"�X<�V�9�8��n��/D��6r?��J��gV8޶�V�T�z������"[lf,�'G�����U�����Խ%jo0k��@��hM�"��Na3��s�o�x����a���1�&�vv.05;{�	o��q�r���Xս�7aByF�\�W/�Z��vv�|�C�(K��ڸGts����Z����0�c����as�}]0g����	�{�@��KM��l���lr�1rx����6��e�r�JL.Ԯ!�PBϩUpxTi�?����_�*B1��_"^���~�2��fO� ��h�~�.�����8�쵺=���V�K�6Oe�%�e���(I�#���t�t�!)��"@W��oN�6��Do�/��J��o�B�,��W��gBKʘ2�Y��<O���/�̓�����Ѭ��� �_[�k|ef��;�o� E��]o��2r���^����y�߁z����kh�~W�}�LwG�݋ɞ�M����^D�9�M����k�_����~Ҏ#+w6�(1ѿ�]����+��d���Q��L�X<��Um�/
w[4(��CR�t�@L���f�.|o��VO�A�6K�IG%\���Df������ck��)_*����4�{���k?���j��NrЏC�%�o:��(�xH}��fX�:��I]�Z���sN޾�:�����������o�LDtW���r���;e控\�wk��X���l���w��l�����$-����v�;�J�BW��!4���H�S5��s~/���vg-(�^eċF@I�6�NfȞ�l�>�>�kd��9����z)�������JEOO�{C�y��ig�6¼���rglt�I�ުZ��n]E:\�3�<�j���6�s��W���I��M�qK�"����e90����W����c\LD��g}���H��=�`O���o����)f���96v�S�ۅ��%�>$��-~�?-5��1��E�$��ޡ�&�8��9���ou2<��U�lݔiH�����cz�=	�K���c���'��d'E�F+�WM7�0*iկt�I�[T3C*��~�	p1���s��v'�_�|�u�:�Y���u�B��T��T�k}���Q�O��:s�����
r��w��)�wf"�^E!�C|�&��B�J� .��.�}\X���tB1�៙��f��W�L��U���*wPki=*�3���q�i��)�rN`m"��3�$^3��X�d�����o��n���<�����x��,h>t���� MT`�W���0%gp|���Ԓ!F��}�ao� Z�^!�Zx�p��-�fM�U�E#(�����˦`����&)��沌�K4�h�,{~d�ϫGߍ������K�m�^NVA3>����D-����Sծ����'y���������([��88h3�h��`@lH�o�k�P�шG�@U�y���k2���U�D �lȓл3��,�!���������ZR�E�-z1�_NT��؎��De���,5�$�����z:�g�z8����į����G��j�'�tuu#�8B��p4G�f1m��ނb5oW���s:Sc�Fm�|�D��эT��^N�Laʣ��H�x��є7�u>eh`�j4� !T񋋨ܢ��%�������C_���)���jC�+�J��z��bk���H$>�wû�➸,Z�x���K.�lV��D�� j���W�BE�6~�e���Ncͧ���Ks8xj"�KՈ�w52�
x�&6���yl�P���ow^�I%X�#�h��ݨ��W�B?�͘m���pOPH��+6�����L�7��[n�Td��)��C�௦���3:���/}�Ĥ�^��!���,7�譀�E�e�#g�̯I���.���S��6���5�c�<K$��0mI9#u�����?C�ȶ�٣�B� �m�����\���Ob�wIȊ���L��+(�dw߱���1���ߝ������0�r�n/{N`��s��r�~afV!E|%0P�L���+�o+$���I}4�mv��9\�J5~jB�vk��q��;�?X���ᩒ9/�ð~H�7�((�6�6w�����W�'�s��	���Iț�?�7�B�T��8���o	}7yҏ�_�qR3 ފ��poC����sΤ1��E�x���8%d��T�Q�[B߈��tW��8e���	]����iS�I�� �Sv��U�Y�$��5��0?T�
I����^��UA��^B���K��׸��R��c��K46��Kw��4��`�+�
��'����튍�8���t��N�4Se{�0���&�^����8�ק\��EBe��0�����,��!����
Ǝ��\B!���&�!�X�4�zw���>�|��3ڬJ��H�-s���g�/���=��}Z1������|Qbb�]�k����ڡ��|���N#��+wr?�
�i�����`��$x@��!�mEg���1�,Q��f�1�dswY��.�an�'\�;b�,Sh�dG5FPL��v���0 ��H	WVV�Z���[5�p�L,L���Q\�'=YIH�����wk�kD�n�<����L�j���C�.ںl���ġ�UvP�Xp�s ˩���qB?��� Ōf���`����6��^S�oꪒ������h�P�\�鿼���;���f��
�s�����}���y�PyѪ�.y�������N�i�+�Mxk��w�<߯j3C<]<��O�p� ���A=��<��ތ12�(���W!����h<d��Ӽ��.�̭�g�?�Hgc҂�ؙ����d垝��K�sʬ����)�rf6!M?/��3|�g�w<쩤�"1Y�̨�!�������@P�ʱ�$��}das�2���Wפ�w�M?E˿ҿ�a:�4�ů�/��L,�����G+�-7�@/�~2�ؒS>�Ǧ������;c�=��Lݓ�. ��"�ܦh�J�A�d}-͔�ʔ�k�yF_�l��DRٺ�G�3������1#vc�� �8��^�6=��8m�.A
�4oY9-����q�_���l~��:���k�� �1�_i�|�/.���"��Ռ�?�c�}���p������_O�x����!�6K��5wqQ�5��<���/)���2$%L+��������ء���L���RM�޸��g)����?>zA����������r��m��KL�c�&<��s)`݆���.��r���6mI	5i�D��4�_���o��x	�bO��ʯ�av��T �	?`�c�?�$K����KD�ۇ�a=���yRm9�7�i,���n��oO7�j��Y-gH�o)K��D&�q����#P�f�?��L���Q����C���}�7��$\��ր�ш���S���,���J��oʸ$�g3�ŏeԌ���}��Ny�����/h�HiU]ޥ�W�Na���`պ��o�3�2���]l�/�6"���V��D����o��z�����Ï'��<�)4l�
n��{H���Ҳ�+nm�^I�?����<>R���}N �
xǧ]e{'в�U�z��ן)M���+kt*�
#�5����� I# *��:�L�m��#��(����)jH��z܆R12�D�-��y Udx�cI�� ���6ZA7�s��\����/�!�p�=Mf+�9h0[2��-��u8�y �AbT>G����Fx!(㾡ߠ�`#`��[�)1�p���̦���-o�ct§`O��YT`��GTM��C棞|�򋷵�0pQ*`t&�65�T�w��I����9��B�����I
=U�;6x3O)�v�����cD&���כ�ұ���5���r�z��l7��s/3�r�J��0�<������������"TC�"'�p6�f����(z�q��m�N�;�-���/�a��W�����I��t�pf�HQh'��*�2��%���"f���;���������q��J�	`,WJG#����RO"s4���"�/H��Yl���8�������("�KbY�{�ۛi����a�����]�|ӆ���ndd��~'�!��D�ˌU[��ޔ�8���8��Z64d]���fH��S�D�����J1P$�`u��5��H ��F" RS9���IQ��.�Q�砬�2�:B��-�ȃ�s���ܾ�K���T��x���+Aw6᲍ݭΘ�!@Ʒ����"Z�}�rM�@�]Z��Y2h���٩A���O<���!�S�d�Ƕ4y��##8g���<j~�f7S������C���5X�Ϟ�Ȳ�ʝ�g ��&w�����N�5�X���lܯv��X0��M��-9�}yԫ���&ɦ���T&Џ���x�î6�	��hۼz��\��T�#"�xҭK���M�gI��p�Ͽ��9��Q++��B!�"��M���|�b��h�*O�J��f��ު}}u��Y�@�M�!##P��]�b@�um���O���DT�FKG��*�VH��|�L�=�نm),:�5l�E.�L�7!��v�������vM�ߩ�c�S@ޜ���-,:�MQ"B$���@�jo����DG� C}��Ϟ=s��.Y�t�ś��ݑ���e��;�O�x~���K��y�x��~"�30�k�e�[�$���(�_�--M*�pH�����e烏7 6�����,v9G\�{H
tJJ�D`�"�W�ؙ����Եy$�;�&=���B���A1���CNa[��"�s��u��}l��2�,�C߻<ȁ�����|�s�>���B�_Bߛ��W�BNr{��Kn��v�zV��`�@�$Ӟ|���90�j�&��F9x�[�D
'I�S��|RS~��N�;p�>kǳ���fj�����lѧy��vl���
��q�G��|m����ǂ��̬%�t0o���۸P�<������p���MyQ�p�^��V��M����pKy��'M1��A��������صq�٘���Om�ޚ���?��b%K��ӆ�U+�d��O���Y������Ŧb3D��L�����FT�3W)���̮o<��c�
���|�K�lh�`����FF���|��26��L˛���'�$P���CRrZ���5�<$��l����^
� >j������
�@FMV�������f##����oU}�?c��˪w��о�A�s鐮4�����BI����F@+��T�z	1Q�>�U��o���z֒����Q߬�iC6�m��(NvT�� ��U����ɴ9�����H�k��W�I��^���8,��m��}X0��F�MNB� &=-�����d�󬏪�yϛ�5����������
NQg��ɰja�`���:��f��,f�̀!�Q�-�q)�'fJ�4o��	�-[���Yb�O �T}o/ i���Ч2���ÞH ��^�o�f5��� ^B̩dҧ�w�^Ǯ��������
��`���!B_B����.x?_��Ĺ��_�'i�_�����Ʃ
v?��]����������q�o3|H��P��2$�|��[kl�iQ9�,�������&J�@U��w̌�Nn��un�-����[<�����x��^'8�����I6��"��V������`6$��0�������G����U��3Q��x&�}B����ǂ�� JbXV=)�i�/F�[��8��7#�cF[e�==@iՁ����u�/z��M�6�PH C�C��p��~{�g�n�`C*�s���$5����͕�`��T�M�wm��Kv���)B��٦ |�$ގŮ�"�S��N&[�:�?_驺g���H��
rssf�YL�ͧhYA&{��+aǊ7�������e��-? ���M!����"�r{f��A�������r�	�"���6CZW�o�7f�!�Owf�)/hz�gQ(�r��{;	@����}Q��8�)-+C �5�*��z��iK E~>(8R�r��3�'����|��M�6�T@���1m2���R��.Z^"*����N��IT���y
*e�\����K2�u������/�4�*�����j|�}M��n��6��Y1T
ȯFR��	~y�a�x+��裢/��biUl?�E��������)�uo[�����Gm"�˟M��O,VV��;z�؏�b?���&�l��^�'
�'{\>�6�f�H8��&�}������F$-�,�	ȏ�����]�S��;�Q�,�.����� bLj�&�۽���L���1"���T���2��0���.���TS���s
��;8���sC��4G]���L�[����ҭ%?�խ�ݩ�h`(
��w>�f��	��TÓ��[ǭ���'{��8��dP�55��C���<���� ����U�Rs¬�ͻ��/FEBI�r�_����P�~�H[#�*&�y��^�{H��6 ~{�{�%�s:V
xN.���߭�X-g�醍N��iܪ�g�T㕁�;��h��xG ��[�UW.}H���߁ر�IϳۢӾ�������ls���V������"�Ņ;&�+OƏZ�o�I/��<�ř��G�r�j)�S�GP~��d��~f֋߂�~c� x|~yy?=�ݭ���-,(�����	�3�2���KVD���.J�����Ӓ����V�l�;�H��1�Y"
+��Yj��OX���uu�B���b�t�����!ֿ[/��Ҟղ=�'�3�>9�0�$�pf�P~_u�T�����񛚇c�N����9��<mQ}��1E�&�V���uboM��gk�-*kg����MQ�� x\sPfq%��ۦg�,L`f�V$g�&�ܴ$��cg�KcQ辪ݒ�C�����}��<�0M�@����v�F�-W&��sc�A�M�����vo���4�@�S"���ʝ�����۟Ar k�2�`?%��.����Y\f�mDLazd~�َ�w��hF���F<�]�)�O͡������Q�Qp�Ic��wnY�w�W#���gC~ȟb$������4݄�0=T2��f��:gb]�h���_h�/yJx�1}�ʹV�(\��7i׾���ѥ����/-/))iW1[*)�4:���Sĵ��ig���N⓸����������}��G&"�+s(Sq��:���`�����]5q,֥���B�i+ݟ�~���)�߮�M"�koW�t��dsT�KF �	�lc���w�"A�����ˏ1��}�Ɇ��z�-��h�!�Ϗ�"���y����A��H�ڏ&gC������F�v�n/�5��W�69.�ǯ�oQY�.B�[q\?�P+d6�)굿����-�;���v��bs1���'X��-�<�,v�������)�g�Y�H�Q����4�B����蝧���6=��O���}��?�O~�a2�WPX&��'C^�S�b����VU�ʏ�+�"yg������2�K�Yg�z
:aP�"����_m?ا2b�r�'(�R���*�f�r'�f>[HPP�X�Ր�����qR�������r��J�Np  �O�#�B2�AQC�S�����P�ϖ[��s��URҜ&x>���}b�gsl�'r�7�y�Ec�IM4*wt����p���kE�G����"y��\B۹60?XK'��t�H�����ة��B,"���	�^�dcB۴U�Gh�+Iw����,������g���l4���a���MQU��-���Q��f�_�~�)�0�䵴�]<؆�g�ZRߎPK��Þf�4u ���Y�\z t��(�g����c	�91e;�x8j����ڭ���.?`[\�(=J��rRy ��q�^j��F*Δ�@J$��rՙ�+�
�Z��ׂ(ORH���-q��+��w:�l�D���D�~���층���0�`]�J�i�VG6�Y�Q�}#[ku��FR���wT|yy�e���A���=>��=tc���[-����~����˦�"5�����G����T��)ξ~~�W�*�ff����aJ+6�����:%�:%_?��z����=oiKPT�M�����o��XN�˓�A5<�u�Jj����E���,''7���}��}f!y��Ԟ���K�'�O23��1��?\�/���Zj��kp�ڥ�b��r�PJ/���p���ۗ,����#	=�f��d����^���!�����-S��j���O�@����>����s9��%�kF֚�f�L����[�d�PlE(���v=t���B� �����i{��s�0�zEG<郮V�Ov�#�Z�6%�פ�7Cm���1��
�ϩ�?0��/3��T�n��=U��>y'-d׼Y�*Ruj*�A������cM�����b�WɈ�( �$T56q��&'�/d���c
W�uzcO��Ч�K���Upb�ׯL�ϹȠw,,���\�5֐Xܠh�&Ƨg�В#�77�D&�9����_ۯ�
���1�{^���e�T�B�o,C���빼�#]Mc����D��"EϮ�~�6�vXPN��
� �����OGp<�����*X���(�r�\��,��¨�s_�����R����k땯���ŗ�KKK�����U��V�����C�M�66�w�?�u���z<�e�{�-b�w��G�uuq����匎��g+Lͼg7��I���A�%�1��	b����2q^n���T.��R3���K�-ǎ�����L]ZZ��:��?���=$@s��!�pe��kcG�]D?���1���6��9�˝��������I����ЫgILc�h=�A�>����1n� ���h˵g_qZf���/��F<��M�>*Z��eq�3)`ڝ�M�@���ƹ����:���;��|?���[R��Å�e�����,x-N���'��k��Q�M;�i�gҧ�>a�HABB�����]�Ԕ�뗠�guC)J�;?�X	G���/ܜ�<��d�+��:Y�R�z�6����p��������4E:%\��x��  f��s�gk��;z� C�*#.��/�]Er1kBi��!�o�&��[���ʅ�I�k�Z�x�̃a~��	���a�2�d�,�Mj�b7�����d�@��O	�����e �F"���V1\��=N��o�bz�E�/�J��{��D$ͧ;ס�/�Q*ϞˋF:î�n�.�b��c���*�������/΋�D�T�%.�uי�[^� \�w�4�q�+/�i���`f��/�49��Na�D�!5��b�&<���,�mHe~m)̀��ڿ�½3����'�wƖe {e˅��ݹ�G�FMԀ�{�7��	ikV��*G���j���b���SE8��e�>�A�uK��5�4Z>m{HϠ ��4�Wċ�5����	9�J�`+�����P��B=�0867���N�[�P�^�
vo��3f�L�5]%i��)���m>^HT4��p����47w��@��C5^?P�^��ş㶢:|c�3�O'M²[?-���g��o}}}	ZE��9��NP�dSII	�Q:�ysl�p�h�H����$����BM05(J�FT�319L�"��Q��>^U:���	N֐q�0e��ƚ�6�E��K/�:�a�xF��@R���3̝��a�X���H��'����L�s�=��⦸IE51)�.��p���ƷC����<��q�E+�eJ+���p�}y i��=�M�.��uN�3�9�r9?�?��rT��SЩU�"Z頳(;�F�*\�j��<߸�=���q�|w~�G~s��8��5ݿs��1Y��㞄dǑ]�6i8M�E�?��2��ňw��v�4�9�S�9�>���)H j+�"�GMO��Y�0�`�h����~�^;ȏ�ZWz��M�Ǿ�Lj�^��(뾤��Ѭ��*G��	�L����m��#t������+Td���Y�Y8�8V��ER�`lQI�4�g�7��!6C�f�o�j@�Xח���
���W��b��XϓO�`G0�b�t�a��e�.DMٳAĜr�+++�'�8�
����O�%�h N�:�F�?IO�%OP�b��j�
ʪ�x?;*���I�j��� ��W�D2���Kdzy4���!�)��IŬq���1�r���� kq���,f�љp���u{۟)Y>����oB����{B��^��[ �A�w��v==�o���ill��*���H-�W�@���8[� �]���F&�r������#�2�+<�S��_�4�Fv���4`�6�t
�j!��9���#�{��_��+a��.��X.�~ᴸ*�������3ҩ�e�pi��=�,�x��B��ژA�ej��2N�_i�(��R��M��1P��㸉��r�=�r��� ���ݮgn�M�YJY�6*d�mK��[��'���;Y��4?�����<��LK:�s@g��il('?�*.¦���6���7kw�BJ��Y�����݆͔gw44�M�0�&R?55�>���p��6�dQP=��e�g��%�&E&7WCX__���O�%UU��L�΍/�FZ�*���?�����W�@�g��t0�ǭϷG�x"��l��.+ߘ��G�ES��(�;ȝ^<����LO���'*�~�Y[����%x<kb���ic�՗��c�fy:dmL�.��)��x�b͕�߿���o��:~�B�z��3��%�_0�'(D��)�
6b<u�Zm�)��,ە��nk[/�9�c�[4��E��i��JOX������s���5���ڤ�4�Q��� � |X\�no!1�s^�C�w���'-�C��k�>�l������pձ��m��R��~b`<����Xud͵��W�i0���L��5Ng����5�E=?�h�V�5�ޱC��W/�,�~7��$�U~\ss>��$QO�|1*�x��2�JD�J2����]�XW���}�͔�'dz���Q��g�Ⓠ���]�fл+JyK���N�&�c�b{?s��\L����w�s�^H��I���p�T��������V�~(��խM���s�4����m�`�y-���P������^#�[/��m �%矁�=2l�lp���'-y�x���w���]/�Fm��w�% ,N�;�Ⱥ�ե�'>����>�=�z���߶�xk]������s�����(K#�H�Ji/uj&u��]�P�dEW0&�ߙ��B�pz'��|7���?��U%Z!:��Ѭ*q�:ؽ/J03�_"��
Z��Y�2��<iA��)&��ڛ��iO����o�,R�q�t�cv"X'��ɴP�py�����I{��g5U/�elT�2<�b2��������0��ppC���v�t4+«���LsG�FU�.�A��q��*kj>���M����3 �F��#ej/TU�[=���z��e�N%���G������RS�DZ g�7a��{!|��p�R�޺�	� ƽi����1���}{[��&�$���pJ��B���C2FG�M�F\��.<��6�rlR�P����\ �����6-�~��VQ�'��O��&�0�,R��Y$�.� ��Q�����	|Y�Ђ5/�x�YB#,���q�MD��Gإ5�t�+}���P���i�������ƕ�uz ��q)
�o{���5�c��qf�n�TgQ�4k+� ��׍��Я"�w�ъ�[�iŤmt��ۅ��B����	tQ�y��!��g� N�U��EY׈� 4qȩ�_�Q��;�ׯ��y���'��ǫ�X�Ť�]�p�;��K&I�;N��ޮ��ωK��o߅�H̶�9��ɛ�F���D�oW]^�O��TEj��,C�?	֌��z�t{��F^6@u��b�jH�H�-���~�pK
����
=6&r{,&�i�X��tꦌ��5l[�,�U�9������v�, �l��K�B;ś1�u�l���MgVzU��W�"x�o����Svе��,�����ͽ�{��&p����2U�C���XO��A�������چQBR��Q��NA�Aah��SJ�N钆A:��.)��n���������pf]�>c���M�5�*Ua�~�p��2#�wJ6��1��,:1�$����
����j�i�}ϣ�A{�n8!��x�J�ۿC���)�CTXXX�v(QktD����腩l~�}�����d�d�Q�:���U
��?���\��e��74��kqc���DFm��a�~��A��",�
P�b�p����/,��k
��\��ٮ- ˲��|�.���2��sV9��|�(�Ӌz�nd�Z�ۤO�c#}/��'���^������f"m���hd��V��s C�}C���sD��)�$<�=�>l�7��(�1~�8~�ȝ��\���ƀˠ�ͫ?q������S�z� tt�!B��2���&Y��Z�������z������G�#F�E,�3n�xe)�w�Yۄ �)��]�B
(LC�����L����I��e��F�+�'�xiv����OmZ��C]����`�v�G�\_v��a�y)��{~O��H�	F^��KS���/]G�l3ª M��%�^���ῥ�n_�Ev���pw�?T���N1�2HǨWR�gv��z�A2��W�bM�$j�~����n��n>�b]�`�a@~��`o���l^ e|a�?D ��Y��1�`��N�8�n� �o��/1v>�Q��.� �>�_�?D�rQ��H;�cK���i*x��G�C�O��7$����j�����6
��(?��\ ���bo�&+"� lD�G��\���֣f��;Q�N��v+H��ijc���$��K��S<;D�>V�����R^�Ƥ ���5��(�p	�����(��ܕS����,6}k������?1%�9��j:�t`2��h���!×��:vuۚ�E��Nc^#q��P����Q#����;��B�_}cn.B��V}��A�
�%�77�l��Ǒ��|��.߾���"����������>-�ã:}�#��x����HrWG�B322�N@	�^�H�\.9��\I�^%~	�0-T�(l����d����8�?�KlőD���[��d��ϼ� ��������Y]�}6���O���D��u3i�`_�j�vM�?)�HHͣ5ƿ�,+32(���3p_��ӊ��V�O�%�+����ܡ������ I^	�(@+�%�;K�K#~�}����9Gʧ\�b5������-eaX��^J�wP���9�鮀=ےW����S��~q�/���킼�CAV�^w$����Mwg\�:��g����'�i�]}��#?m�s��']�N^:Bۘ�5.�w=�7�� U��X�������"|�QbW�.�׼���wp��4<<�1����I���&�
?7�"����U"�U�t��́�p|bj:T��A<)Sx�Y��c/�4��Y�.]屫Ӹ㵐��G�X�s�]5��'�`����wz��},��n�|)#D#��J�%�ġ�X���������>R�W�N�Y^!ۭ�U�b�z��H*��s}�O��i��[^����k����s2r����p���*U6d�����g��ݎ�_�W;6̴,�J��h�zNj��y���&>����`�u���!wiZ����f�߳1�i��اy�\��4����))K�����:	�K���kR.�@�>�����js���K>����x�JD�"���R�����M"����!u!�����^� #�����l��2���Kp�Q��mX��;)��xn{:�����Z�%W�B�	<�����}��?�1<O뚂�bk�&p�@���/��eCJ#�]*��<�A��p�P���Р�!��ɰŕY��M*K0�W"��7#c2:�l��ڬ�6�}C�OX���^�.'��ه\��5:��CbJ9)L*|}}b��h�C���j�N�R,����y�^���e��ʆ�c��k�9�X	 M|g��
nu���y�����A�?l�Q�^��\Y2u������=6��ʑXܑE������vw}3[G���U���\�ZR\�9�j��Ď��_����`v�do�h�NV��:P\\R�Yri��~�V8,�Xh�7H�T/�w���د��(l)a�h�Q�s!:k�-�fe�A��yV��
�B�))����9� s���H&Qթ��3M��g�B��/�R���Xt������!�j�d"��	�N2S|b{<����&{c\j*3���ij8@���	�A��TP��r��$���Ez7w�N��+�6�9+�TP�7`�x���ޅ�U�#uvv6�R��U�^���ڲ�aV���q�������O�L�
����&����Y��;dz�����O�(&��Imgn��Nt�C	q;Ġ���xmt;70�ۖ�D|�)�|�d+�;��c�75mk����[[X	���с<in|!S�k��;{�}�|k��h�aq��\�PrU����Q#BG3��3Mʞ�"2p�J�j��L�%OS�uJ�c����vb�E}8�:����4G��22н�I8i7���R�57GS-V퇅�C5����+�Lcޝ1���jG������海Eb�^���|��(�*�Qu��E?+c���y�u>Ͱ���ߐ�ޒv��sVF��E);�v��*���.���p>H^7l����t/+!zD�G�l}���Q�2>
��a�cz�oKf�-���N޶��׽j���.��z�����a����m�or�\��LyB�VP!��ۿnF%Ir�/�����;���C2%.���\s�ejCq�޳9�j�3����-��B8;`y/�>��6�M�T���������蠹{I�+}����J�CԊd::�KS�,r�WQm��lgY�k�;h(7\�}�ޏ*�3j�M���8�8���$�i���,:j��Y;<j�2K�KB�"?8��xHR.�,�(���yO,�h�+�����g=}*E��\�rA �	���_j/�Ş����QS�j�5b�]���4��/}7��>V�p_s��D���2��4�@}!I|� �Q#ǱUR��_]g��=�E�&.�v��$�=�׷�������.�il|e��y	�b.����u�D�N��9��x�6vϯ�4���rrr�RR��N��c��T༛@>��0?S�>܈'�)���p���V��̜5���:��켏K��
�"mU�Ǒs�avz��f���=��=?�낣W���6$�E�孛ە�K�ҳ&�N��z�\�&�.�:���}��T��)��-�iN����#�|A����k�N+Z��3���ǰ���;.S���G�8��$����q�6<��L�[����p�t2�>��|rQQ�S77�)g����T��c����4K�ٔP�	4��4L�as�+#�@�К���r+����7�D| 5����6]�r�SZ��)�M�l<=u���68��6ihZ���[�:x�O��ZB.a>�Ɍ!x�ū�UF�?�Wχ+Y�z|q'.�u<(z�्MJJ*�v)�n[辤�xȬVX002��ly5�w�u �,j���'ʴ��I���� ��_<��^��&�sY8&�K6�S
����ċ���l��I8m-�$*�n�!�@��-���
L�����"�_�fM������P���.�/��D�AP�E8�);e���!D��5�9�n����7�Qÿ��F��8A��\w��k��Ri��#����Ś��)[�B�T+Q\&Sab+壼��e��ι�n���w�B���v��s�ۿv+}����?Џ@,�WF��}3�b<��ϛlq����6��8��g�$��Qj�h2r��Q�Y�P!�BXճ" j%�XG��8*�� r�̂[���j8����}��W��P�{�P��ޖ2`�A�7��L<�o���I�,��w�aN7a�v�7�˝=g���(Uݶ�����y=ޤ�7h(y�MF�$�Fx�Q7�z0q�Cq$��5�w�&��4<�J������]�b��3�#�]i�ۡ���Ն�G�/`������(��3Ieī���<���^��q��h�\ӭ��/���+����_{}��2��)��}C��E��ݍ��0_Z�a�4��y�\Y�X����L�N�UTT����V�'rx�Ƽ�O��!u�	�<�
B%Ǘ���>�kǒzt�� ʧ��IbX;`NZ �ą��MɅ{����2-�GU��g>��ʒ#�(�]Y}�.����L�%$sPS
�|p�ԐD� �M�e���/���ĂJⳀ;S'�>�9�� �P��}���ǵsm� 'ܕ/�+%��3�+۔41jy�O-�7$e�N����y���%�E�S�g���C�	�����@3tA�}��͍6͞�|����A�~$F���(:T�d�e�L|��M����	m��i�^��?��ݹSGQ�!S��g3�:������X���.hO�o�p�[c1سu����WL\�8Yʢ���b�?�	ND�Ql>�:jX��
q��?���%����#�W)���W^�i�w�P�WZ
�d�5���J|�ŭ�QB�� .~8	���A���6��D�M�Zc�ޔ�Lx�vґ�6S�&�_0F�+1d4�q����,�	u�P��}��� ��5-M�6m�7Lk��1%,b�w�'���3���zF�^��L���&V?��ץ�ｦ����=4��m��N���I�����g�������ܐ��UF8z�-���V�E�Xi�	IU[��M��;;�5F��۞��QĶ���ok}��������.�b{�,9����{�v���,�%�Dh�^��ib����CӸ�3������$ciy�6���P*����O��t�[\��������<(���D��m������h�ֹvy ���<�Se�594�4X���C�Dͤ���,�)HT���Iw���}`5Q�?�=B�U	j|�/f���^��q�A�Sl��p7+�_�4;-id٬)G�
"}�A+<{� ~��as^�������8��ͅo��6ܦ�c��G��BW��7�}�J�_J��8o�+ ��,��r0[.P�t��Γ���v�J��(�S��PoZ��"�F�Ϟ��\-�w5��E���F�C�� �':��A������W+&�i����F�bO7L3���*����i��,����>�޽�s��UZ��I�n��[j�ZS�CU�H�	nR�����(X�/��X�k�f!��j��m}R{~�Ph����2�,ږ�!��PvU�*�OG�*Q1l��s�N+�I�������r�$g\h�sYVq�?�@qb�aA�D��ʝcn�|�f�W[�gV$$!]������V�{�Uqw�����]���w�!�c� ����p}�Zlw��锠\� ,hN��4Zt���V�n�'�W�}�	�U�-j����o�t9�1!3X@�
#a��1ٖ�;]�Š�b,�u��z�/�Ď�fA�?~���˽�O_�9f/"�0!zC�C�����j�X�`��O��ڇ��u�,w�]2���j�a�����<:��Yu�ygNa����),���FcxW���{+����jl^�xk�2��ޚ���@�U�umi5
E�gQ>�K���uH4:̯}�-�>�S�m��r���@E���C�zuj�:q�\܉MLA·�9�j��\�=1)���V�
"��<��«K=������L�g#��10��ph9'�.F(�@u4 Fh��Ghhe?Q6��<�����y8�T�5�`�o�|�/Rd�������hz����{������o�+?�a��RBF� �$�k����j%�w�"?�� J4)w���ͥ������g8��l��k�S
'� ��^���W����}O�'��~X7a.5����������脓(��P�Hdhoω�_.�7!0�D�w�jWB��kB���F�ӱ)�����xyq�Ț��<~�Jo��
��	�8G��<�9��oT���7�����:�YC~SD� �����B����m������Lۘ�_�x�@u���Ńm,�˻���!��s��LV����j�c�o��P�cC��`����W�V���n�y�����@��ނ�8%�Q��l�U��j�E�Ǜ�	á�i7�2k//��p������7Y������^��iȲy��Џ��t��:U���}����H(�n=n¿ ���]S�:�%��0>4�/���7i�Wx�TR��뭾�x��K�"���f#
v��_3<Ű������H�!)s���Y\Z���dڀ�|x��y쐼?zz�b�%e[���0�ipg=�����W|�:)魤��M�vl{&5�֡�G�*ax��&�(p�ٓܨ��6��-��/O����N�e��x ���vJ	��{�5���q���"d�æ�mh����k���}�G�������uE5+�Ϯ@N��ЙF�?�8���SA2�X��ɘ6�|�7�Z��!6���g��j~:~f�޸>׵�j�FΏ_�Gӵ�6�r�@<������b��\׾�������R��" P���8<'.���0yC[<��:n�B�/��O�zc�1f;\E�aq�|DrP���j��*DϏ�s��.#L�~DF�;�+]�����j��פd� �3n�ՅøLos?l5�C��5���hnM  ��-�t�oG�x4פ���=^PR=��H�/S�3z�!��*�޴�����;#-�A����^���Ō����\|��¤����`�P��`0�ө�����~�@��3�I#��<�7'��jAɹ��a�d�]z`��� �+a�و���OC�#���vy��fV,w�e�%(i����&*���rz��:C�h'�12r傿�{@�����XJ�~�Vd�h��4#�j��iW�s`VCN[H�K�{<��\��Q��TfV��]�m^��όc��lF�!�9ل NF�5��ԧU��~/Q��������ʱҴ�.��|Rz���5z1�k�����'Y�7o�"�R=�����|_�4��^�+�!i2\��I�����p.9fW�&ط����DOb>��ǓXq�zzH�&��	4x�d������1e�K@M<�E�p�x2utgw�;Ԕ��/�x�5���Cq�{q��`6%^�(�2̜.[���t�ƴ��էO�+��,ر"�b��U����fy������6E�O�����[�9�8����~��}!)��$�M~���hnc�q�v�L4�����p����q�D����Nh�1Ud`ꯧ[py��6Z�� s���m�J������=�����>����6�ΛՃxOˎ�t�+������ҫ�#��ڠ�Ј��w��x<d�DHn��i��g��o+g��m9b���nm���4�����Q,�iba�\�SV	寰��Jb���0���e�zx�+����"8"�M7�5�����s�W6C˽���%P��Ύ��|�9ʸ�����T/����E��=��`�6Ϭ9�
�8 {`��_dAA��Ke���;F��,Ow˅ee�lӯ���I�{v�fFSK+�ʁx�d`�z��}�LM��~�So}���]�l�\�p��C�gW��?�_m�0�}�y舌~�pZ�@������^�^����T�4C�:[P�e�ih��M���݁f�M�ZZ&��X�k]wdQ;����d��4Ѣ��}�͝�ͷF@N���������J�u�l``g҉�ߥ��Pbv������z�� Ը�Y^��Ϋ+��_=���~|{žv�3N�C+�Fڂ�����Q���Ғ��"̎��-n���9�|x���|��H������3x��n�-��*�����T���i���_��D-��w���{5F�=4�4��ض���kT���������Y�6-fU5��9��ן�=o��d�u�4F�!Л~�kH���O����m>�p��-8+��\dl/ʔ�J�~�o/���CԟZm�s�_<�1��0��yZEM^��:�c? �����K�I!�u��#���LRix)��qI��*x��j�T���O^������ȏ���)��u�~u�i����v�d�f[zQ0���q3��v傄"�d��Y��<.���qR�|A[F^7b�?~�D���{�l.7e����t~�?[=�H�O�)�.��,���r?8��^t�p?��;V�{/�4s!`BѰ�j���V"�U��GbQ���k�%o�Y���B�}%a�O7q��Y38�ٗ�qv	\�v������f0�{���ЋY���<�D�b�>GJ�6�������������S<�F*�"��ݝh_�-�x���x����a�5�h��"��`n�Mr�'�MV�c/���^��@��)�6 {Xx��^I�On=6ru���;lY�l}� \�)y����K����<w���)�s�ۘ�-�������}�A�yۢ/���ꂮT�p��x�9�L��@wJ ��d��}�)#n��4�ڃS��=�:�X����r���k����ύ뎁aa�BKo`�~������7d���:eDj=ss�L۲S��BQ��-n�ku㒙��^�s�]�c&�E^W!)S퀽�y�s�5&�'�""w�Ko0��*�$ܑ?���lʴ���mtd���j�Kf��p1���Z}_i�M\Je�w]XX�=�7�J�R��)2I7r��&�;k���H���h�x�'��i~D�[Z�j!����B��F�[� �D�w��e	�'��(�e�jO��6*��+���N��8 Q�&�a��&Ҧ��{ۣ�;��p�u������ԷX�����v������G(�n\�݇��C���k�ϓ��=J�.J�Z��2���d�.bS�b�'����춱��3���k{�v��}ԶY$�$EJc�K7/����N��I�Gu�?���#���R�%
edj�u���㪓��>��ڥmo`���[�ι�B�o����Fq\���T�z�p�t ���Ti�&�7o�u��䄅�9�\[��]���e�ˇ��o��q��nH2�ݎ��܅��f�b��I��C$:�6=!)z�9�s�d��?�܆�W�ܤh%�|����R�Ϳ�.%�R[ØU�����yf�0j������e��j�a�"؋{��}��,膂�` y3���n}m��<����{T�@K�ׯ�5�tb��r��yJ@B^f(1/���B?�Z
�w�V_{r$a׵״ԕ�i�|������a>���Vg�OKN.��G���=%���.>>���J~���ᡴ�Lkk�x0�_AU83�l�O���f���Y]�PXQ��^w~�|@#>^N��#l�����s����3���\L�T+�Hw��z���?���?
�!*���.V����z~d�Sc��9��oOM!�ܬL����vK�P�~Ů�4ZW2�H��jE[ß#虀��ݷ_�T��^H{�l`����k.��_-��"�����|�|y�����<1e�jz`Of�ɮ��,�ͻ	����zv0pߒ6E?��?�P�*���~����~xk����h0�0h ]�s�}��s��ޒ#W�cJ�I���#X��g���R���X�����2Q�
?3�;��pw�#}4&�&3>����sa33���}�"��������Ea2���Uo����l|�Ƃ.��jĊ�@�vG*Ed�os�9�څ�l����d�^p ���g��B���m%o���LZ"�R��u�W~!9�����=����v�Ff�1�So�i7��+�0��6��k����d�W�_*A�i0��O��Nv4羿'm�Ub-\D�Ծ����K�mZy��/ ,�_Td��bj�fxb ��B���^1���Q�h���-XL�%7�)�1��i�������8�l���OOh�\{ ��Sw���ysǀ����Q����gZ^�{��xMT<�<	�-6��'I�;X<��~��\�TY�Mg��Yͨ�J�%�l� �p���$�����)�o������]��D��eK(l���)�&���I���o�L�z}}���	1	��'*�;v��Cܾ��P&�,�9���8�8?}��+U��MF����H��3/�~��f|�&�X�lB@f{�;���;�G�A X��~A����m�).�Źs1:�_c����������ak�ɽ���[�r�\�H�O�}�8�k����ST�a�t�G/]���ĕX�~V�&@g&e��C,�Ȉ�{�Ģ+-Z�|��:W�SW�A?Y�w�J%u����r�G;>��{I�s&8j���jK��&q����ή@��6v�f6f���i|u�mykF�,<(ê�]�4��?�o� ��G�}���gW�Y�I����d.N��:7��:낈�%��`���Q��e%���Tt	.m�z0�Ƃ��ʸ��]旴��G�BJ�I^�����<�޲��mص2-	@?�+��� ���|�{2�|u�>)&
M�`���g�:L}k����-�#�f����k�O�r<�H-��7�Ğ� lU)������TQ
8%�z�x��t�gR���{��}r�4�+KĔ��k�7�$Q�/>�Қ��9W�告����~�UC�	{$��L�%=��ߙ��.��M��Գ���Q����U�@ݙ;:����a���T���B=���n�����.K���[{��nb��Ζ8�� /5�7�8g'��_Zc�L��.#X.6$��XV�Gɽ����?['U�
n:̫.1���q�(q�ynz���Tc�����!���R�ѯ4��	w��:�P�L�:w�(<�U��\!��/�R���P K�G���!an��C�XCJv�I���k���E~e9���B/uǸ��yM?��L�	pq�\Z�aJs�u-C��j�N�1�C��b�M�6K.�Ő�O���Zc�5l�)�T�œ;]��P�D{�y�y5�2w�W�Az��گ��pF/ʜ�X����@����E��u2X~�}ł���h7����IfM��7��<�/G��6$�
E����<y�~��%�׹g�<��/&���#���X�i�!Z�BJ �Ęť��߰�r)�-�뿅t>`Gↁֻ���1^ab�����K�	���|l,���7tŸb�k3؋�F����س4��G���=<�'�OK��ūR��Ox��rP���ǝr�g�{��;<m�k�����ȶg߾"jG29/Қ�I7a�r1b�ݜ����ZN�Ҫ��ޓ��\vm����),��nR�/q@qd��4H�	�f'�z�'F\���TX�q�2oy�����JZA!�
����ի�H���W����/��r�'J+���C��RcH(�u�K[<e!ca��e۞����ãǱFsΗ�-�Ce����q��+��p����5��u��u�8�w��l�����o:d�_�<��y����4�W5p%*3�\�7聍�w/�|�g�άύ��xq}}�����N@'Ͱ- �8zaƓ?�����~Hn,5���!XcY��aW˸H��-���b:15,wŭsE�}|?�),'�*v�w��	K�����Ǖ�l���T$��dq�2�~�VV��ONK_''��uz�X_�*:����a�m!?#�z�q3���5���G��q��k��6�Ć���I1��O��$��G�`Ii�?3P�����_mX��&���F�?�bG{����"u��N��@r��q�!h��������f�r��G,< �=�g��ma�3�a�B�;�J$�z�^������\��=Kr/x���>a ����xo�}��*^��٭'���ڔ(��G2���"����&0}�a�i���x�4�[�3�f���_�7w+�P�>x[S=y�
�7�گ<�!˃�i�n����F��$\0%�&%2����ª܂ZG���g�$��p%��cVI5{ ��+g�1m���#
�O3pYUFXW�Ͼ�=�X��4���{�чxZ�ƒ�hƭzh�I�es�&�l����ݠW���^�N�2J��)Lw�+��K��r������_�]�W�`�;O���-�3U��~4��X��b�M�f���bm��BR�<�[9g�L��r�/˂������MQ���r4�ť����J�}k���o/����õ�vi��?	�� �2C<t��a�j&��~Á��-�d�kݗ!E�<􄆪��d9m������+*�:��V>�����Y�Щ�Tϑ��9hd�7@q-��7Y/��_-�Xr�Z��]:,GFb��b��oS�\r�Vf��v��p�x(��c�r����JC�o��/9Efݻ�������yy��#���7������^o��L�w'�O��"�T���*�G����
�C�'��F��B�b,j�|:�#N]3#�ĵ����=��ψmӯ6��\��X�kt�I�9�~���(5�N7a?{9DuЗ�lX�TY0&��	~��Ux��ֽ7&�0C6�UY��Wܼ��6O[#dd�����	�rZ(_7k�ÝD�;n;���K)��B ��6�[=Eg�h��	��3Ew�o�o�Q$�d�#��v��g���/�����B��̀��z"���d*����5��r�O���Ar��>�h��n�����+znY��[LJ䕺x�*�/��HW�!M+;C��w��y"��@vl9�+�Z�]t���,��:�i�t�T��%hT�ц����<޻t�T0Y
�H�-��\�8�$I/��j�l1K�����'�.�8�8D1>���޳��~>�`hb��;�'�៉w*���Q�30:�#�P���
��p5�Θ�/]0��p�:C`M�����2���v	��ω}����)U��nR�Q�&����T}2Q�ր�X�%�� A����k:O9F�[�d��$�-�u������7x�a�O���l��t���	����E��'��}p>�+�SA�-Q	���:�Q��{���gn[�OD9e�4�@N�-��7����l�r&���݃��q�_�����Nm5���)QzR�z���q��v����%��Ǖkq�Ŗ���u�����Y�Ý���mW;8|�Uk�r?`J/����t�5�!��9�A��=R���jϾ�8�c�ӗ�;s~p:��V�M+;[�����Q�4�5�>�͑�d�ؘ�����BLOW�a�z����r�eѣ�a�����;�B���/�_Ƴ8���|��K�`�a�p+��C5�D�n,9ԋV�����6"E7� �� �|W�e8c��\�F��-�Q��T��&,4ڗ���F�n2׶�w���Dqd��cߺܟ��u�L��90S�w0_׮���e`ް?c>_�2��$��FL�ۺ���I4����a�/���{}UB���$�.\�B�B�vm.4b�nUd7�A�w����In^���p�c�4/#&����LLM�s�*��+m�0VQݡ�b�l�{�y#p�����U&kN���Z.[��+h�&��P�KK �Bհ|��[`�r_�[^>� ��13[\�G�����3�5�qB��������^�x�|���0��z�98�X:�RE�,0b0t�����+;<^ݞ������Q�%mW�A���=�a�+��&ey�T�pL��uj�m�t�]����`F �������ʠ-�_-AE����I���!��ꝫG��k���َ�%p5��9��6��'
��{8��{u�����)�^�TNӰ��Y�݋��:	1�ޚ*9~\��8�8)Ҹԓx*��ah&T20xv��o��l.�ײr�����`od8�����ug~75a5a�~��^5[�#h���Vk�C�p������8M����ұ���`c����z-"��-�)+b��Q��H�	py��A�ok�:6_B�8],>�l�<W���Z�5}��7n�u�(��**�Y�S
�̚��sܗ�G^B�}CVL��&@f:I�Š�#�� �w����Q_��P-�-�D�v>��Bι�h�vx��FZ´v��J���w��9����!q�N1����d�ɖm�6��{l���}������/����^n�Q}�4�����+�M���ye%^|8I��	[��.J˳C5����fdD|Ik���dTdJ�J�E��~c�g�$�rHZ|I=O�@%���ճ��`����d�u={���Õ���k:K���w<7G]��FK�Xx�L�b#w^iLJMH���G,�x�(�/��3���jLC`�Tv�ElAS=K,XA%me�۩w[�ɇ󉊮�/�Y�ŦG��%�yg��@�������vP��ᡗ"�i��Ɩ�f�Y�! �u�Yd;ē� �;�]py��~UN�]�F�n���MM"H$�@�C��|��L��
'�}4��V�������ʯmeQ�7,x$���kYٝ_�J�%,�(yI���|�Da��;�x�G���Y;�$~"�. \��7�#�=��J�'�]㧷���G�ͦ�q7��R�O�n��|j���C�ƣE�dq�\���'�������O.�rum�I���첞��T���"�Ăr��H�$rթ��Y�!����I��V$2
���G��T�YOʸE��w`��h�=X�-��հ��Ų7����ql��0�T(s��q%#���>����[\�M{����>��Q�6��<Ii	p��7&
��[nh\c
[nk�����^!�~��s��J�MN���� �!�&����R���u���	��T�_8=�:^�\����i�a�S�=�MG�N�����ݫ�w����Y�M��<�vO�x���}=�������!�*6*
��g'ڰ�����$�ʶ�sz�}���_��	���(�J�._�ז��~+vCn�z��_�D��Bj�2|+rA]�ƃ�Z�r�N@�>OaG��H����`F�'D�cV��zv\6T��E���t�ms~F�t�=DI9x�ۘ�Y;��1�l�vh���l���D�:�#su�D���,������Z�*�	���X�e�T��l����'����ԑnCp��U�~��WF�_��6ˌ->&�M��/[�,pi*--�U���Ը	L��\lm0=��t(�Դ>L�b�Ӹ��&){�O����6u�>X�SXޔ��������?�S8�tf�S<e��������@�3�ג?)�ѝ��o6	=y����x�'�����ϧk|���'���C"��##;��qSMyyy��1W��6�e�Sl�6�1|׬c.*���:����-�D,�t��> .�����S���'��5̜]���d��x���c�u5���+��Ë��EI��~n&k�X�k/~��Q9�6�3�F���M��T{���ԤGC�]�^Z�r�;~�Rܣ�ǐ���_7�aċ�X�j��S7na�Mvwy�w|�s�>�[�����Ebff�����őL�&)�շ5� ��f�<h	��,&`��Y9��=���x~y��-�y��^F�y!J�:���>(7<r*���H��������d0% ��,�pC���P�F/�f��+��a��z_��&pP��U�qY�I�/��������J����c4�93a~�}�Ō;8���;�p�/z�M�&�uч^�������>����{AsːG)�y��۷m��x*�**.{bZ::�#0����q�rL�] _^�_�6�_��ډ���T����ߊ��qb&��g��W��F2��k�#R�h����?��8�E��y�i^�L6�BlA�y�<�}�K�[�Z�ƨ2�'�pE�Y�^탆�	��y��J�?m��ף�OXG��^�F�6C��ֳzEEA!a ��>�J����9��i��PkO�AрU�UT���(#.#�Zw˙��%G4R��y#G01�"n�b�?h3�Jɰ�v;�ִ��=֍�.3�G������i=�x݋v�=>��ݶRv&�2`��g�}⫧]����F�8�J�u;J��$�.��2=-2)�g9V֩u�3����GI����L�o�\�8�u�I��.����\��m��M���g~w��d�E%d��dڀ)�M%����t> �S�l�������@,#
NdŸ���v<�d*�qQ��M#���-k��Wd\��O&�/���<.Z"RW�����F��� �W][��Wx���e$H'�T
�s����#�v%c�pct���=|��`�����Wƃ}'�y>t����,���n��b�o�ESc�d�|�M�z&�oii�Kw�=a%9�Û"~{(����K���(ْ��]{a�G^�ˌ��ͅGhC-��@��ˌ}Ï�`^��^���H�N�O�>���9�l�qC!��~'����"��;:Q�zW�r�ܼ�#�����E����K#b�`D�'Q�����Vx��Шk�Q�N�������H�;�r��4|�a�#pB�xE+�����o�*�<���_���⋷^�������XT�/�;{���R0��D����\�k�T�E,����s���:�L��YƯv���m�8������ѧ(���$+% ��;�CڹSr?��mo�G􄰲�6?�߭Ơʾea�'|���>��[�q#o�+���no�)R��O�~,� 7�A}���ea������o9���3����MO�����bPt��B����}�3�؉Ա��5ރ�9�$���u�CZ֒���e��q�t�=z���}�UQ��/�8j��G�|^�C������7�^d����I��JN7_P! RT���$����$�L��Ҹo��\)K�������6R�y9yK���֗��4�Y�3Q	ɹy�kV�T�eX�[�?L#!��(��t#��ݍt��t#  -�1RCH���R��!�0�������</x�u1{�����Z�0z����D�	0g��S��xTN/��sO���_���%��_mcJԑ���X�N�a��ٲ��HhX2��I��@�) �)}[�AFۭ��kvf.!���Cf��ٮ\��t���ɗޚ gL��&u��Z�q��,\�����mi�B�>��Ij�H-�(�<�rF�Z��aj[�Tڗ�D�S��;�F<F��I���Gp6a�A)NO~oV�����Z�t��Ѳ��>�vP���;!��)}���Ǡ�A��D�cǏ�;��0���%����WrC�����$��X�xM#P���ޑ��m��0�+Y��g�`M�}���-6���H�B��}A���.�)�.�1µ���$�>Z����%e���%���BA�丂^�T����
"�yo��YܢN�<���rÔ&�O��s��{�fS�}F8� �$-&ZD(���M��蝄j+%�w��N�#���I�l���0>���Z��=�(�_s��~ �d��2�C#��sh��?�T+b��_q���Bl�r�I))6�}7�K&��=AZ:	S|�!�6�" ؝lO����V���Nm*�F��P"�����D�xla�naI���Z_2��D��CJf�}�6�/M2={��h+���P��wgdA�jY��{tV������S�\_�ם$�[_Κ�]LⲆ�����ҫ{����Aǫ���Vm�R�{�%
�n��w�w4�������b��wM�L�h�8�g��"M�8�ӠT�	�*�v߹�UZ�<Cn�uy��wa��B�{���Il��т�q���6��Zoy~)������/:ӊ ��w��X���dX(�}�w>?
�Γ xq�����uH*�P$6�B��tR׹�v�*S_�����I�D�>�����R���3��r%�6Ɲ�@�KS���"������ə���-�k�P#<<>p���ycEVX�#>��pk2ʤ��L~�Qo4^�v��� �����ʬbt���²�`)��N�Cx�kvO�lcy��@�k0	�C��Vt�H=v\���CK=�0v�jJ0���k��+��	ӂ��2ؘ�~�D!�n4#��6��;&!\vĈd�!gp��#V(�h�5��0���Hz��'B3�+r�F_��>9������� ��-Δ�W�����ǅ	��N���������	�p�f[��&�T�;�_~�x��;���3j'�������Lac�U�ͼ�}N �+mϏu͖��A����Rm3�B܄*�Ǎe¹�e�o717?�>�_����c����C
@V�K��|D#S�̌��J���3��`��._�W폞-����nX��D���'���\�n��bͻ�?��5�?�[.*h�t��֖-odK�)�%-�:lJ�6��Ĵ���4�g�薪L�I<��}�B�A��s^�Zk�zE�C���0��/~�p�z�V�*��n�S��¬�J�Q�����Ќ��!�p����ö���5�4�%5~F�.ܧ��ݏ���ܰ/�+����ݜuRSU3hi��B�v���ym!~��Cu�X6���'n����6iPϽg,|�E+�WZy9C��f�<��x�0nQģ[;__��Kf�������&��Ć88��&��`�D�6����5�ܰ���Ү�������h�p+������1`��[ʡ��MwY�SK8�G�xKZ��J���	Ji��oC��Xp܀ ���#�2^�t��V��[3Z|m��NҠ�d�(T �z�;���;d����h����שWֵ	0:U�5��o�����KzLo[N/�5F�`棵����E���Gy��y���E�'&����0/�U�_�	���޿�:T���,a�L┽:-Ҷ�HIK#u�hE��8>Ͻ�@_� ��GT}P@ �2{**��b��'����/����&#�a��6�ؓ�:��tP�ն���U_�x�6N?f%���hXz�bL�\ŷk��bǁ���T�˷��f��������ߛ5�����pt�$�_J;l'_��%E⓾l|w�x�&z}+�;4�s�\ƿ��=ƛ_myR��P����T��?ko9�~
�ǎ�b{S���FE�Ђ�f�JKK�W���`���}]g(��'����A&�{��י�i؀��d����:�1��:V�2��S�Db�d�	��v�[(yg��J
�t-���'���wD���Z2��|":��>�����Qg��6*d[�'�Hg��PS��O�^Ćap��� Y��b�^K�䷟d�Eք������VA��e��G}��O%%��4y����?$�g5��Veى����gi���t>Q�cTQU;�Hb�� ��-'㐤���|*$B�/��<��e���d$RL!E�I=���pe6�wR@ޑ��a�p���[��
}�$��o����5k��@���_��Q�p���0{�*�Q"aH-{-�T�K�=K�#�����%z^uj}��u�����ЖE,���3dqc/)�^�Q�7�;��߉���������.���N:��^�f�G BO;X����]��./�v�h��soP����'�;��lo�d��:��$	qh�y��L�	����?H�o�ۑ6��x��Rc��ǃ���G>=gq	-��{��A����ނ�[jē� �T�ӣ6�����q�J�FX��ף��fU:���?��w�sr$��]��d�B���J9R�?�x�k����`+�������ǌW��`�j�Q��a�Ɣ�Y���[��8J�O�� ކ]��ԢR���7E����~2+�������I�Nr��O~u���O��ێS��IQ�[�E!fs��<�㎊���H3){��&�����L���x��܉��>�	$}�����O�1D�ͨ�IU���zW��{�����2u��]O3��u.I.Þ��+�KPH^͸�q������8�Je�9e�d�����j�[��Z]�ͯzS^��g�F-:���U�X�a����Sfp����
=AYٔ	7COp��W�d,JJ���r�T��8����:�WFc\���sr��oz�MY;?��L���{��u�7��+��L�3�C��G�<����寒򵎣�� ���w�Y������w{�)�GK���R�D� 8_`�c��Q�o[��r)8��M@�3�������»���� t� 7���1�������fB���Q�����@x�0�߳��|.�,hL�`���ME�B�	P��{w���V�j�t�X�j�c6�[�?|��֍\�H9�Vs=�	�	���BM/���큖�;h?`81VaTZW��M����T��.�ݒD(��0�盰�N���X�>R�Ѱ��-�6U3�b�@�*R=e�<���~]���05��wFvw\k��2�5k��V�L$��~@7����j�]�y������Y��������"�66X�&���MV+�u�L�2��k�Q��"�6vv�����@(�e?Q	��񉐭��J���fS2$�eÝU����p�����q��k0���	ц]�����<1E��{n�	��Z��AP�s{� �L=�b���rW�<��~����>/�u�3о;9���3.�:^�d�$��+�9��!*��4�Iԫa#�k<����7��j0��R�:C����7�}�X�FF�$���f���.a0?�Z�W��
Y&��3/���jQ�KR��'�Mq�~1�}Y�`'�OX��Py`������2��/EC���W#������@VG�5y{�j��[<��}4yQ,+�_��L�;˦*���{(7e�hODc�R	���P"�O�!�|+`�7h��o�w�!=���.s�4vǄ�!ò��(��OL��2Ѯ{.a���R}���fy;2ݴ��e��[��l_��b ������D)/�e6�e��zT���آe%���q@Q���I�f�WQ��?ߵǔ���r���$%���9�k��V�d�w !߻�)@�����~���U����m���o���fgz��7��3��Z���"qta�RR��I###t�H����~U����'!)����������{�)>&�᝹:c�FN|2y�3p�z06	����"����B1̒y|��*�H�}���o�X�d���6��Ï˥��Wo�zuT{we���<����d��gJ:Q��'�/�"^�kf�N�v�c�+~���|*����^<l����v���.���m����dz1��Oѳ�'���]V�,�\���U��J��$�W3��5��3E��dOP���x�sV)�Ϥ$0;�yn�(C!�Yp�WN�t��=
*8|u�<픤o� �y�:��Ȩwa_�!^,�׉kp� ������ry�8��%�5�
���\:t�����R)Ļ�~�&�bT�L�V�"��_^h]d袞�Iv�S��B��Z_�2��#�>א01�mX�k���g�=+�<�p,��E;��@��w�����¸�/����I�O����k:�H�!�xZɀ��|�@�\SQ �lmm%db-�������|��\X ���f[�Fyr������#��V?�Lv�@o��������݆��a�{JL�tFz� ��Lg[�'����NN���M/��k��2�b�7t�h����,�E��S6��Z]����<klP�>v{�8`��=��O�E}rp�n�_�S��{�j����J�/B�iUu5؇��p$@�m-���I�)+v�=�X��Z�'�0O2s8���D�K���ۓ�m$�*�����F��O_z�O��\�Q��DI �* "�4H ��qɳy?^���]!C����py�uǽ���%߰^!QɄ��[[�)��ɓ�I�����Z����~5��4G�j3,��t�t�Y��O�F+������㟭k��cSS����a�p[q?��D3����+��Zfe�+�Z�fD�w6�s�`�a�[z<#�:�����
o��G�_�����G��#�Q�a�m�b'����%#�F�1�]*�)����A��'�!����0�����`۹)�����������7�!����]���*\h�U�)A�ɻ/e����l/�׫�����@<?#EUE�9�jaar�yy2�� --X�P�Z__���.�.��Kk����{�臾��x(|A��6�B���e��{���Ĥ���-!���G&��m/�_E���u��;�c`q�LM=�j��	�L����� K�/�n����S�s�ڔ����O��7�*$�j�!d��	�w���aL��'��,����C���O��c	5eN�R��D+��-�3%u��WM�\�8�F:�)z�zwjy1<����U)�U��9�o�����~a�{���y#��y�=�~�'����s��w��d�2V�9Lw���^Q $L-T����]���L�j�vޭ9)��^�P�Y;R^=
���:l���z������I��ex^75���~�Jb���������<0�E��O��{��꥚���ib\������;*�g,��\���ed +X����.�5�r�W������G�6��������/�R�G��~ɮ_�sx����0���d��r�@�6g���0b�h9����c`*�],��0�����3t]��#{w�'Gb����;��-k[eb#�4����\�A���gE�x��%�j��N\�������RM!f��&@��7�<�$pK��b��-�@xM�`V�0���r���崸�R�SO�1���y+o{��)K�����O�%�Nm�+E�3\dW�kΖ�i�=���=�n
��9d��R�i�jJ�r��Na�4��U���"4�#DN��9�#�krr=Fee�#�9NAA�Q��`Gb��L��ш4;<$d��#@�	���b	�}�����e���1�g2�)T�L��HRRk;'��r�Zh�0��<<2���9﫩����㽰;\ � pѦzu7��{m8����w�I0��_Ow6�=ǎ�/�l��F��F2M��p��^�ojf�^����mc�� 	���ڈ��F ��Xr����!��Px�/^�m�;�r�ca ^�� �<a�,���f�m��+ٴ��b�yMW>�xM{��N��HĐ$Y�O+��ɜ5��T���	�.~��S<t�%퍤���}����6_xmooW��3�AX�Ɔ��V�i>[y����v��7<|<Ai����7�4�h���Oϲp��jK��@��u���!;+�/f�/9������=��oE���>��ND!66�c�`pYX�-����.©�T��[@G\�d��S:F���}]����U�%2�5��W�:�`+�w/[ـ_�
'��G2�I�����͕�V�F�%b�Svo�agD$!a�0l����ޗ�L�z�$
��<\�{���!mԩ�F�93��|����T8�V{��C�]/��?۰�T���Q��B�LYYa��+�B�jy����T����M�G�	�#��֝��Zm��p�9�#�>G�wn��a,r�bs�X!#�=>�)�m@��c����%��B�����a� ���>�����)7��3���n�潕�k<�6���]+ߦ��O�Z��55�8�)Ē�l2��P��m7mG7��Z�Q�ЅfGRIIɲ��ψ�'E\D;�,b7��F���u��5fTy�^ASJ[
���]cϢą����5�9 �׭[�ݲE�g�)>dgZO��V�s=s~��_L�T�����w�K��R1=^DMB�1` ա��:SZ���S%%�|ji�z'�ak�U��}}F��el��;�"�D�/SI�~�-�������,���KD�j�}���
�ʕ��5�x���qy�O&�	k �v���g#��ԯvK�0O߻g���x��(Tl�U.O��W��c<{�����ASzG;Q�8�Jdo�}}�=���3��W����>��� T7���f�&`Q�/�]��"���8T�* {�E���Gc�f�z�CO/�>xv��/��8�{�ZUt�Ҍ&{:4:�ibb�>�TY����|Y���6*���-O�p�wm+;;��EC.�����45[UU�< ��yx��%��Dd�\��" l��E˙oqs3��R�M�K�E��pB��qo����s<tr6gz*���=�{����Nm.��W�L
#�Ap�D�1��&�H������㚏�1�gQ�p���Y���W����ܾ�Tl<C5�}�
�ׯ�(ʍ��C}�GU�|v���ztG�]f���i\O0�"���6�`�KLW�Qn�βC�綌sn��M!O,\�JDWk��R�S&��-�7��>hu�=�[�Y��&�ޯt�ȷ��ҺNgf���X1�s[J=[j5/̆� a�0���� ;�Y<X��8��ώ����T��B�;+T�[�`�-â�&6Z�"gqf�>������a�������Y�p��� R"ù+5c����c8�&A.�C8��Y�_��+�<�M�!�����@�p?�d)��.��v���������"N����j"�]�⌊���;;���I��|��ݩ������h���SWG����5`��Ğ:/|���	�;�k��#�3�(_@��B�@�u�����Lx��nq,y?��ο=(��6��iJ4�0�dp�.��Gk��\Ȇ����,ߣ���ӗ�o�L�n�Ok_�/[��4$ y�0�NǃZ�xR�������ӊ�f�.'!�{V������Kl������W�+�3��T�;/�魥X(�s7�yl����������ؖ�ص���,���n�w~2��U�����cXHt���
���Bd]uף� ���p�h�D�_B�V��m3[����OԎ�Q��������X��{�7�r�����i$����=Q������D�Ǜ�+D�f���;�lV�L�
m�D:xV'2�V�W���WC�����{�w���eb�/�������,y�0O��1h�Dʟy�(o��C��M���S����p�0��nQU�!pR�3f�8$?S �Y���_+�nIlf�o��B�"|5c(���_'o�aJ嶚8�N�9ԏ:@>2���(�鷰�8�z�����[m�7}�cr%=��k����Ӣk|II)F]�!d,���w�+�at�M�s�.2��5���VN` <t�pi��soមk[0����߫���ҧ�_�/1Z�����K
�X�����!�@~zs;Y�]Jŝ�#G��������i��C ��TTT����WR�'
���D����k+|&��L��f���M�ϵ�8�ͯ�04�Z�����l�m�x�M�l�/��^fe������;�e�\ާ�;}���z���i��zB���?�O��z O��Wi!�i�}V�c�8V]九-�1�_'i�Lj}CA��!�;� �}]%ů�\�Y�=3��9��n�j����Q]�*�����G�}�F9C��q }���T.AF�'ȃyڃ�p�_�F'���O׮���Y�r-�vҠ|�3z��&,%������J[3�IVN�8��b�ޱHh}��n��dG�u�7�+}h'`&��հ���SA��c�R#������Z�@\�&�g��F�c�[;lv�Uƾ�_ 4(�B�oY&����F�:��ޖ6�ܖ7E�܇:�M=9�ȏ���`�GL���T�9tI)��M.����w&���F���nM�u����x���gAPWbA�e�3_�d[�t\��O�c0�y��ɬ��T���g�j�M���Z�P�������Y������X�`kW����Ŵ=��v�^�9�z���u�l�R�^ژ�����%�U҈��d�#�q���n,��oP��G��ƍ�����j���Eg�n�<aŕ� y����c� `���v,���2����&���{.K�E��q��'F���2��8L> �p'*8LqN���1�*5g_Î���<��}[���
����,��=x��1P�&eb���[y������`{H���ac#L7����'��饈>����.�XTi���Sצg96yz�ƓP���[Խ�>o֯{�`pi_�#
��j�����\ScRXt��6�s�=���$۾�f�8j��SƸľe3�F��Η�S�Ь���"q%�?�@yE��b�B5 4O���IBϥ�Y��刯`����{���U���� �F���t���/l�J�قf�^��s��2�L]��H����/o�t��|-���(L������дq�^��4�U�?J�gy*�μ�}`�W�|5zKmcbc�Ng�ĩ��) {���p�r�i^��:�=��9� ��IJ�ZQ=lԩ�<��>�pʯ1'�b���x1TSF�O�3��)��}�kОM�����R�?��'/t�r��7Ęo���S\�ש ��E{�ԯ~
{�����w�@���G�2��N8X�:X�"���'6vKO~���U�۝�d�^�����)�.�d4�o��/��ܖ��'�^0bE��e�[��fl�!H���7�ӏ�[���z:n5��7M��H�r�vk��;�����{��� 'Veoo�����a�_O%&|�9- ({�;��^�v<*��{�Z�
S=����ݓ)���n,������Y�ۻO|"���AE�WB!ɇ�h��#��w���c�ںl_Ӻ�m�R׶��@?�ig��%G�X��U�pG����ZK���#+?~Q��S.� ���AS q9.dH�����H���ݛ�o���|���@p�,I�{)O�?DN���8�I�ox_8�0�=w7G�eevoM���wM�x7>�W�<�=�Y�������b��'�grl�,2(�3��::����c"��:<�yF�C���o�0]�!ߟ�\��	=���!6G�/�rFq��Oh�Z���a��TG��g9sT���[��9��Ɍ��*�rm�tC&��z�[���a`����	�q�Q�P��)���|�k��{�p�6�tg�z�����+�`>pw}�
�z��gNO�z-A����>��HtTvR-�n�� �j���Ĥ���:���m�ٖH�~��8(���'Se
R��Fz�e(-ZR[$�YP��`T�I%�u3P>Uu�2,��xb�_P$��\���U�A�N}����&�/�>�a�Y	:*��Yy����kۛG���(�¼������۷��JY]�l�9��h�|f��&��Y6�2�wq�8���ĚK�"\&���ߩ�^�������=*�u��N�E]�E�@�����ͽ%>'�FVo|�U�{��o/m<ݲ�_�Ϩl@|�2#��yĊ�v�N��!���:���O�Nt�4���Z�\����wkFB�Н���=�;�t�C���E�C�����������:mtz�Ɖ{���mh'���C�\7��Aq��wؐ�������;5���y�\D�?G�kQ!�޻Ab�6���j, t4U5	�(h���_���	�pHߺ�1����	��Խj�b8r����+z2�GEA�p�H����s�Xs]��}�gR�mPG��m��s�n�B�������ϟ�m���9�op��$.�y����ָ坠L4�Fx�e9X�F�hq�ӈ��vɴL7%�v�/Ci�� �~>�-:t�^d�Q�HS��[ʑݧ������_��B�8��i����Ȍp�黿��^`���N�4�VR��U�#ď���8<�)+�vIe�O}=�q��8,���A��#�#��V`וM�xH+#����A�R��z����y��L�Ċ��]4x�9��ږ���uG�E�ތVg�7��8���$ r�螯?{'��6�|;[�cP.��(��h��/�j�oku��
d�T�}����m�����3���I/M�{Tz��)�?� ��3�Q�-�Ɵ�A2���i�
� z��)����PMOg��&I�a[/��_��g�|[,������p�.6!�Ch���x ���D�`����B��cߧ��'s!O�{[kʩ�:ɞ�=/	\���vJ�����M��}b����z���ug@?�NB�ރi!�ߖ�U���<g���v:���/�m�݌I&�u��充[|��0)�4��(�~LП%Ŏ5��F&?DxG
Lo������].{p���V���WٟxcX�j�ƝTQ��b� �П�X3%�V �3�8�&<Zk�D�,���l�uT�{rd�DY�� {V������2���|N]�k8�u�(*��[#�����zqj�&��a2�y����isr��W���Ϗ)P�1e�U�����g/w�?����LR��(���2d�����C��_2�Q��T0J	w�h¼������~�x�v=24�r��EC{�����w.��{�P��������+�$���Y���ӎgY�:>��ue��¶1՛1�"�^���%\~Ad"�7]#�ȭ(���	1��~ݴ;�
�ZI����5��]E� ��]'6_X�AY�=�|U0��d��:���݀��i5O2��O���[NE�ZY*8׎��/�:��a�
����WЀ������[�z�O�SLI�w�}B����c44vx닐r2/�Z	5�*�^R)~����~�����R�=�G)q���o����{���=*$��_5i"�7�-%goܗ����lr�KN�����Z ȗ����t6M&���) Dǰ�U8ER�-�`�ߠ��񫷟o�m�g�Q�2ӳ���8C@�AA�@
z��H(s�Q�W0Ц��	He�� ű��BU$�Z֚��U@���_<���p{�(���N�ޅ�CKwO3�G*�1W5���A�&E�������)�������kL>�D�,5&��z�{�-6�^�>YC2�w���,�×[eP�mfoǢ�
1Bd��:��?���~L�OKVnؤ�U�E]���܃m+s�0��L�<�����3&�7�i������Ͼ�x^����j�&k]���|��>$h�+y~мS�qp*����T�@�m0:JЇ��2���[��)�kM~���B���yG�M���M#�����B���(٭-�ɋb�e-U?�{%���V��\�.=;��m�����2~�T��~<��L$�g\8���Z^�69L�M��c�B�I�]#��!m#�σ��)3_����vE�lk����q8س��jV{�\ʱ2��+��x�.��������K{�Iar�ĝA��B��1���l�_H�+�ф�곲^=1b�`�c��_������6� ��/X>�V��Uv��-o�x"4����4���&)3n��(d��B�z5�>s�za-�n���&gq?<�yI ���ɳ�#W�H}v��p�V��i�W�_}���99��n������tϭ�I�{�~��t%+{P�u�V/M�t��4��w�������S�ᢹ��b�4,�S��^����n7�鵫�R!��?��M�|���Jm�Rf06���{C�s�4iD��=d�6�|�sص�T|f�Yh�ޒf��K�+ف��|�{�O5ܡ"�?uv.�߼>h7��p�Jr8�Q���<��$����i�7���_��J�E�ռ��c<�	Y��V�H?6��5� 4|�$s��X� U��#W
�)c_t��8I"vū� ��G�XM�쇮Qoh��\k	���;��Q�.���@��.d�2�߯l3���e�����UkM3*F˸����`��wΥ]@����G��;����o�Lw�������v�k�I!�1���;ˊ\�hS��j��<,�R�p�N�e��Ƈ��˖R�0��!��}��Q$��[���Z�y��ҭ�8�r}����0��mʤ�@y�Q�/Q� ���q��c;�)�9>b�gP����މq��
C�l~��d���d�i�6��W�=����m��c���Ο>|f��ܬ����_���7��kDav�)ᵅ���g��BBdzN���h�ke#�7����m�\c����F)��g��WU�(�'��:��+;@4��QK>�[^�d�Ur'�l,�N���mp9iߗ�c!�^lc���E:��D0u��@<eS!j�o�0L� h̀c��_91���	w\��  ��Y�H��z='�ZH��n��|Oh�`nr�yr��^�nHҐ����W��*^A`O�l�Ƕ,�pCyEMQ ���~��5�կ~�Q\��[� <!^��a�y��|y��)�b.�.-��"?���%�e���z��� 5���V;{~*8���
FBW[��S=@�3J'���U�	��}��YZ����0w��l$t�y�q�b�>�B�@��X��+�m��}]T��M)X��K���r���h��|���Q���{��g<�ʝ
�k��A�>7��)QN�V&�ט��>�N���C%%�)sn��wk+|чK|�jٔ��f.�J[�ЎUe0��a�������>n�q"���pws�Py;vwE;<2�-��ϟ�^_�ȩv�F���e�O,�~�������#�ͲX(4*����k�"�@���������f7Ə�K %�G��jumF�/���3��/;s�Hŝ:N����|,�/��E�s���~�?�����ō���L�4l4���L�Vq��t%��P�q��W:`�x[q��.�&~dY��yՔϚ/IL��5��T�x �"}��/^�����.y�%�fZ�s\�Hp %�	�>,��Z�yk���ׅ��2�4ǡ�|�?"({>  +a�=q��H������P��zJCf"�nj[�5;�;?�J(�m��ƫS������?1�#�
�#����`��+��G~��5|!2����x�r��Tɱ��tƍ
\8���lw��R�͢���є���m��DVN
G�;�kg��q�	�s��\/E'�(�q�RΦ=��7Mr~]+G���?J[T%�7n��{��$�3e͐>�k�q����7��b�2����iW�]�(�⠳\�m" ɗ����߹�7Z���F� �+j�(l��c��j��L0Nxt�4�`��o4q�ڦ>�¬�q)l@D@�FqM�zA֚���(�\��eG:�{վ��30��Tx�{_p���wE���X�*(q�kW󽅳cU�r���ٿ�
Mʞ��*��	NF��`������F������dd���n����eP����w�S��߁@GQ��:UW�����������)	�Z���x5%bfG4�5A�!8CeN�~��?�z���υ궊2P��;F՛�7��vN�����<�����L��I[^q��tKATv{���'[�iF�i�,YF���`Sח�ɏv&���rOt�X?��aLa�t]*d�l0Zv�W��A�A�L�L�`��:ڤ(P��~nE�v��1;�&6���J��r"
�`n�T.�u�}�k&Ch>�*�k��e�U;+EqS�Ǐ".B��2?d !BN?�;V����2y���W���U��>���q6�qy�1���<�\�0�n�aLaWgv�q����9�����.}]!����\}r��)ͣ���=��j����R��	�V(=f<�k�fA�n��Ι.�U�D]^C$)$��o��{_MlL�dwJ8h���F�jia�mu�j���Z�2��>����F��^`�9rPӇ]����*�
�1]B�a�������Lj��f�:AI��ON$��6}m�&d��
�u�*s������cb� Qo�t�����R��$�f(��Aa���o�j�+M5�*�oh�U�g6��jk��qZM�?�f�O���M�������'�F�s�Y7͵�8�_����jܶ�V�G���ݡQ@����������h�6���>���6�={�u}2�2�K�U&�����bE��F2�%�.�-W�I�Y��dDK[�֭��1u��r�u��Q��և�||:c��/py䵚�ij��=���+�A���]'	��2��#�krX������e�_���-����u�,!m���(���(�����!R�aYki�kly�'ü}bT�������c��7u�'��D��	�ix%��+�Sk��&� )�f�&�*(&%�F?k^�HD&�Y3B�qtys �e1���|n����®�����o�1��+��;ٗjj�{X�c�⟏0\���)^�T�̗/� ����rW����Q�D�$�n����}���m����D֋��O���k������X6�����(g���<�����l�]?���4��O�X�k˶
��0����E��q������?Ǫ��C^L�엔����FU-H���y��thp�?9�W���.��B�>o�qb��������j@�f�p�]A�� DC�����`���x���ync�z6������y�4��_.ڔ���{6��a�8"Q�L��#��/#��Q�I`
��g/��������<q�I������������^�a7~f/�g<�Pƽh�=��-������T/&����u��z}�C��J��'��?�+���#��o�JT>e������m�R�r�[�}U]MU�i7���U떕d�&S�����C|���~�T�]Џ�?	���)�r�7�4x1��������~QD�yB��i3+�fd)��C�;�	�݀E��,i` �s���{i��7��?[je$<S���cY�`U�׿��*׿��c��9��*{�aV�.!0J�g#�L�V��c:�G�**\��(^o��(�հ�US�J��I� uoE>�	�F� ��f����ui�h���o�q"ZחE�h��ZK�΢+��&�������T�-⫔�1k�K��S������>��78�lvll��'�ITܔ�u���}���TK�fvl�HE@Q5��d	5
o�d����5�kQ�֔�Rq&`)��mT������ݗ��u��w�{��J�q�7R��A����X�7%�� Zz�������2��8o�ɻ�]C}j Ǌߋa�hqF%$$Ե�+<
����i_�wIGU�\�!^ғ�M�
{�~0��uB��඗+����T��a����$L/g�3�a��X��� FھokZ�N�n�K�A���$J�v\�n�l�� ��KGf����{��2=�S6t4���u��Ń6>܈2��t���~�<IBdtt��،ŏ%;$|����a��'#{k�@JW�C���غ��?  � �a�Aʹ�R�1YEPX �����K�6|��A�f�\�G��J�����:<�.@��-^KpY�%oou�]ng�&�����w'v�ݿ�'�U�ї�CA��?�[�/%��.�f��^amc߯�oŋ�ABT����15%_>2	�3��`�h\x������/��;^͓������ZJ=#��\��8NK��`oio�h�F��y�+�8Ō2{��"5Z_�(%������}�d�;H �ʞQj�M�;�4���n�Q_����a7��~��|�3��Ia���\���ݻ��Y~�^��✻��W�UWa�ə#�\�ee {zz�V�n�>����G�)����i6P��	@���T~m�BP���ؾ�u���2+`#n Aw{��;���ш_�$2�W��+��X��!毷V/��uK�*q��jެ��費-���.5Yc�0JF��-{1B�
��=|EIIY�o������@�:Y�U�<�Ƣ�m0�2����CL�Cp�mlR����>௦!<�����y�=+Ǵ�QE���zd�� c���:�=��9_�������G*�H}���q��������L]��͹���l�|���z�k��~\���¯�uݒ>׏�;��S������M��ׅۢj�ޔZ5kojU�Q#j����U�gѢZ��,�v��{� �.�D����}�?�~����9��s�9J=_
��q^q!Gf���*Z�_~��W)�CѺ_�-�&$$+�ᨊ�<��i.��8Ǵ�����xs����E{���G�Ը�{,�Խ6y�T�D�W7d圣KA�/���[Q�@��P!��b�Dv�|��~Eyu5"����ۯP��ײ��~����K���Ŵ����觸$6��½(�5��pu-Wп;0<� ap����ϧ��e�Lbu�v���ͺ���e���v���X�#pBh�zlNWق,����O�|�G8
�G�9����Rc7����X�4���uz��Qg��8L�:��*��N����p��PG껕�3Û?ĎX�i��f�"K?���m�J��cLzx}�t��G���2�q��L�-��7�_�PG�����x���0�~-,Th������\���SSs�{'`w����b��aT��b>J*����0g̕�>�es�zaR��#�t'a3�j��N$i���T�mG��>�l�yZ.�� $��z�*�����s�2A�#˕){�X��9]��͘��d�[OHO������AU\�ԁ�I�e�v�<$����2?�����9G�A���R�:��+-$�^�X��������7t��N�v�./���!gڰG_>��>RF\�}�.Q�u��Ӣ�><�&�����a4��f�����KV�l}�TCBҶ"�la�.(�nڤ��%+�n,�~{
[�=^7a)D��L���%?���;}�s���yHQ{E�D"7.��lc�T劌����=4�E4����ަ��>m�F $�n-P� ��c��!�b���r�������)�g��d��~�������踮gl�Z�"h�iQ'R�Iԭ�Z�
H
�g�	��ҥ������7���_�/E��͊��\Fl1%�O�Uf���gS6I��[CZ��}je9.�S�����J-�P��ƛ.�(:L;��E��J:����*�X��^��x�5���Zb�e`U2�l)���T�봸����c����O���/`�:�z�I��������c=B橨����(����g�Wxڟ�$�/H�gK���ݘ�Urjm�L���#gu
��m_��[?��|��[!hZ=NNi1zq��|X72����"y�*���K|��@\�t��?T1��	�s0ӝ���3��'f/2�}g�ZI��K�2�/C�V�"r���d���#l�d����P홍��Y��lgL	���ψI1t^��z]�^zeQ��,!�j����(�k�a�,V|��˨����Q]
� �N��C���*����S�D�����	���s�Z��}��ɟD)jG������S�&�}qs����y��3�
�.���'�A4h����`�j[�k����±`�E��M$�d.�R�����x��B랉S��Fe|+z�����lڂ:E�`�X �qa��g�&�/;���~"/Y����P��{�w�8��fk��yB^N�z����������u��Ie����^���D�����?��66��L�sb꭭n�c�ЪZ�oEd#8+��oڭ��;(��&H̀�;��O�T��
`Ig�2�#J����H��Z� ܰ��:��%������[��z��L|�#��ϫ�N���%D��{�y��jIF����1����oEzb#�l��:�6q���>\�_��`���ߋLD���nC��uk��0�O��.J|�U)J;#n��:��8Զs
���r'ӑ'�/{To�iڐ|���������!���xGT�秠��)~o�DV[���}W��߈�k���1�����sttD1���E^��3��X��y��X�=Lc{�K	��Cvs����#�輻�3;���j2�>k�����`|h���Y2s����KT��+��ȂuJ�4-�[��$Ҍ\j�r��O]�]d�w���!�XVyZlEf���'\��L=��;�q���.cOg���������Oš���.�-��̜-`�"�b�8b�C���q���C�4�B���8;Z���;��f�烼WG)�+�ߋ��L�o�� �<h�{�Iԅ
����cS'w°t�:�N�tu�@j����xsj^<R����D?��� ���W��Y�c����o�'u��
b:ְ���C����۫ߥ�)̷Ǳ)���ψ<�޼���WYƔG��C|��:/�|���U1��[�������8G�z�����o���F���C �J܍�]�
r����F�����k�>��
���'�*��-�J���\&���<��OM?,�38u�e��]E�z�o<j���q�<cˤ��<{Y�]��y���������
l�<���#z�̼b�.�*�x�p�����,�|rK:���:r��]2�+ɓ���K�|@@������S��X���co��j�9�.s��r�)�-�ފ�12������6�a�>������ǫ�v����^֓���K5KtV�������}�pY��?��	���_��y �w�ܤ��.4��{�Zyؔ��ύ0�+��	�<���jĥ42�X����8e�$��ڕ�n�?�l�-%[���֗��I���g.aN�C�_Z��J�Ը;�b1�x<�O�j�e������(�]~ki���WQRz��[�)`��q$S)k)d��|���!gD�0o<]�dwߒ����f���&иf�ēBpڂ�{d���o��U������"���=@�}	��T���=
�s�a0.�)���Ϭ�E(�CNc	�2�ٵ�}���?���:t�DəC����nm�K�<F���0�Y�$ä4��#W?	;H��T$&Yi�_`���'<k/ŗo
"�_0�x��@��<`Y�e/�7G�B��;�/�̷#F���j.Y2h�������6�W͏���ql�k�3�"ޚ��*�)n=�hf�����mI�}ڷ�I ��~���t��������O���������b>N6�֮Yhz�9��vY��9�"�6���7S�'���b�K��C��Ta��魍��=�q����J��h��A�?�5��X�z�,�BH/�^�qD���q�c������C�^�U��Wm���|]�4PGl �hF8����n耒}�i�Lo���G�=4�6ؘ��I��lnT��oG�d��4�oE|LA��Ӵ���.�i��2��(M���ֺGQ4��Ҡ(�eyRo~5a�?˿���0^��\n�+HJwW��_R�Z9`"2ob/���$y
9,�,2~��OnO�m�X��PY����7��Xg�RR7-�n5|���-��_hp�"Y.������L��IQ	()�?s$
M+iL.�_]@���Z�֬Q��u�>%.��4-]���&:(��T�6��T��xY='�S���OP���{�7�ǥ��vV����j8���97t/�hyς*��8��5�m�h�����E4��d���c��h�ѹV|*����G
�w!�$�͗�Õ�{���YX�Vp��&�
�pe-�PDs0p������O6cIp D�R.�(dN��i� ����J�����*S�����!-��䬸1�x�f$��@�mP�<j����%`%(e3}so���������d��<^[�S�N�q�(�:�`N�E�� /�T���/Q#�Fd��G��vա�_K!��T}i�bџ���������ة�y'�
�~r����d5�%��e��F|z^&u����Y����@�ި������YKk�i�6?͙q�x�]�/^S�`��0[
L�/�����* SS�¡�����%^՛6�\F����͗�1�CÂ�(ɦ������%���O�\0�v�A�R�����ӿtc�S1U��P�o���&�r��(PF��*>i�շ��!ۘO���+
�9��ח����
:$�mM�̡���_&��-$`R�f��k]7j_�\�5Ñ1�g������R��[	�gۥ�q	V��ϡYq�!H�9؟P%��2y�Y���~ȺY��OW�vX�xBG��|-T�tY�;���G�l�q��O$�թ��l���Ӝ�l��C{���'�ԢeK�9���f�
x��OAa��Ѝ���)�/X ���4�?H�eJ�r��������� b�#�9��A�[mW>w+1E��u��;��g^�
�q�\��{9����������|���M�' ƛ̈́�u��񞰣Q�^Y���c�b)�Dě�p��E�9ju�GsE�=�B�S~��Wى\�l������m�Հ�HG�In��,!k�f�b�#�v�cӒ}�� m��ju {Vw]z�/qu�NN��&����ZE��O�?���� v��-�k�mC|Y����[�G儙�e
m�f�+��� ��X�N�$������I^A�ӊ76JJX���'�������~�`��G|+�DC�8n��8����Ֆܦ�,N��秒��M�Mw�(�������=�3��-��g{���{��ʞ��bhʤFj�y����r4��obAhf���/��ux]��(�����<Js�]}�2�WQ2r���`#�a�HK���-�^�Z\dpԽS��k�?1�
2ϫ���lu���a���v	6#�C�{���3w֚�Tª�}�j��4�.E5�u��y^� ~FjlĎh�L��n�ΞI" ��,�^�ǥ�]n��d-6�F�~�$����xX�=�^e�dI![4k�3�&(#���πIv�8�Q��:�)->��T�-�Z�h�d{ZFq��T�M����J���je--"��Kk�OB%l����u�N��`�s�$��YKy���Jz��j�R�S�WU���TQ�)��9�S�ߊ��H�3�����f�P��IS~����"	��h��@�o�|�u�_کljj�h)`=�Y�w�}���^��|
 	�^�|G�ȍ}�݌��m�z��]>�D$�����\�СN�ͪ����'_�q�?y�vE䓁DV�6���K��vYHk�ݗl�"'��+	���hgE<%H�F��p�a��}/���ɷY��7��-���������V�����e�����w�{����������M/��?z���j�{;���¯K���&ce����[����s���)�+T��G5�� ռ/<�8���u�T�a�U���g��5=�zWQ��s��Z�9�XH���΃�z�\	�=�\q#��it�^��=a�H��_H�j�1���n�s��(�2��O���B��i3���iT$n��G��л�hʟ8Dl�l�sq/���.���t�U!}ι/.�M�|���2��L�R1���6$b]��vN��Aǅ��S|�4�� ���
�� �=���H���v���[���b̕���1����~^Q���N> p��F6!�x���җ�:�L�r��ԟGȽ�ԩ�R3�� �`��8 �0�nz��;��6@�Z)��NR�m;QNf��~,�ޖ��ھ�dY_x��B���sDD=��W�5�t��D`�u=��I���;_�E	�,���ܚHk�8���ӗ�/�4Z�ih���齌'G�.��PH-.���M~���]hl*z�_s�]kR����O�ݞ�>�L�#�I�k&�-+#b
�}�����Cٔp�5eZ?k����5�׆{��[C{���i-�ʶ���as׷���V����kYJBε(��g�J�DFPo  G/=<jꙋ[��=a�.!���H���;E+��=�WKL��٣����Bo���Vu"��nq)�4t,)L�#Q]W(��ks�8��Ӹ���z���i�2��&�4 �e�E"@�ϝ^T��y�#7���D�<;���ˮ�Q�`;���K�`3l�^��<��̉Y^�s�w���A��k��%_�=�a +��o��%<��Wh/���LE�����
>�o�xE{4�t'h��1/��Z����R!���LY�
<��_4&����2{O�y���x���+��Wl���G[�d����kA����$�]UX�+�%���^��H&��D_��E�Ć9��2�E��qHcu�]��xT�"hY�i���s�ՀvL�It����f`jʟ�r��5|�uN.[�����.!0���Gy�ܡ+вE���A�����;,�!�^�7e�b
yI0em�]5����qU���E/��Iy�R�t|�{̣A��pW8Q~tt� 3�{+!�T�0Ǚ-ݯ	W^�G���<�0\A1_���/��1��})��eNqFb��9���jo��
���p���#:oKO-}���>��76�-8G��͹� ������w�$�
by��L�]݆��g<M����A��o�4E�)S�q�&2bx9	�y����w���0&0�3`X�r�u���H�V L������U�֔�9��)$�6��qSKKIL ¯���C�ʵꯛ������� �@^Ycy^��9��F���Nq}@�_�ܹ,�	ڽ�x�����K}�r��;���qdFF�Ѽ�����( �*�aYZ�$�|�G���%��j����#��'�(�<�O������yq���N*�%hմ�[`�n�番���|�y����G��¡�ЕX�omr��������OH�=WH��v�d������aA��aQ<l�Op�N^zn����n<1����2�?.���|�!�C��N�gi.�m�XF2O�
���+��Z�xA/H��s��҇������v��Q�^��=�5���r�g;c�*���o�	���X����~+���P���C0�-x�@"�籶�͟WD�	^hu0�^w�kV�M*!0c@k� Z���������S�(�q9>�UͿg�Q��O�M��(��cm���.�wy������F5?��`���|�f� �,<�� 6՚:�=�'�2hn��'B��[9�$tRy�NW!��t���8�:�|B����` �^,Qߐ�;����ѣ�F����3��]��ʡ��C��D��c䈙�[�톿u��xA�#ALK�;��Ñu:�à\�Q�N�����j��U�P�g��a��;crON�d��K,+^�,���p�b����.n�z
f��I��E�y����a�U;8!�N�H�o9�����X��ёF�w1��Å^c�Pe�Cg��G���R�^�����n`�L{��!3Z��P����K��lT?HU��^Z-�Z�E(���wg�Y��@Ҝf+�����A���0OBQ�
`RI��2G�����n<��R��G[Ӵ��6��>�c���
3���R)�%�
��C��J݇�R�3����'o\S����0�-?:fw{�q�ס6s�ς[A�,~�K�����NN�!鎓7�L=p�4�"Z�j�A&�˟A�/���fW1�4�v�O��]�d�<���ݧ���xm:���9��^o~�X����*l����,K��v�z�`4������H�j_��`��\����#���m��Z����r����@�,[�PD�S������G�O�/�.+�䀤{��@�j�^�iW�N��n�MY�UN�Eƣ��'����|�m;9�A�c���q��d�ۆ������^mx�V���4b��'��O/��O<�������x��<�n>�]t�L���<�Z��G��-��j���S��_m�x����W�^��E�t<�'���ł4Bz�z�-Ɗ���~Pы��}�P�!1sO��-h����վ�WA����wz�xk9ˋ5����-��
��=���2#�r:�H� ��C�SȎΘ]w��c�$�T�����-����2b�#�O�_I�d�Ҡ,�O0Ζ��;/סLb�ō~���~Do7��x�R�ٸ4	�ͩ�0	И�!k/xD�Rb{��Ίm 3U�E>۶H5�Gm~����9@i��G���� u�͋�� �����侂
�_ BA��ohƜ��.�9P�v���B���a!���h��E4-w<	6�����F�V/�r:�?{x�Z>�a�t4��Bs�c�%e�*ww}����y�*>�C���YsJ��?�\9�5��"���ʺ���姀�]���7T��w���?�s��`2���U���V7Hhf��<�VΘ�:�����!�n:��^��n�Np��9c.���Ϸ1 �2�X0�7�7�Ь�XJ�}�Q�Y5�χ��[�T�jܥ����U����_�ks��k�?C��pDGWF�5�T�*���[�!eF�0T��{����� L�����ހHDkd��u�s���s�o�PbQ%C�2�}��O�����/��,.XHc�+��������_�p�z����70rR>�W��I��p��p�/�C�3ه�)2Qv�f~�9�ɭ��#���83�2�
��3~��D/N�*s��e
�����a�/h��@T���mg���wڄ%X߹������(@��L��`�5B�z�%	���KG�E�|�$q[F,vZFCdF&H����l߅ �;7=�l�\/T ��PЎQ	�{m��@JV�w��"G�p�ۮ��]Z��j|�W��ъ'��m (��]�G;H��2����D$hj�>����Eܗ=����+�/L<f�ct��T�D�GlW�ѕA����ס���Ն��!��E�&_lKF�u|G��8j�|˖X�Zt��&yGE�Q�G���yB�n���l�@�nބ��O�[v�hP+�E��)�I�D���a�g譂G�=S�xE�}�&�H3��J%�O��*���]��\k�Y�o��6np&͟@�\?*L�&�)8���E�RG����a�2X�>/(��2:�	)��|G>o3;	z���8�KlvF?�A�T�k���/���jI܏�]���x��p�׼Z3����U��<�M|#�~�mV�.��	{`�쮊�iӇh!K9�����y�X���%�Ϛ��+�1g�5!%2�,S��s�Kd�_c_��>OHK�:6����`v����|�h�F�e}�����}�횙88�"q����zw���Gd����g��	!�p�"��w��"��@k�(��p�m�=::�=j�'"�^�M<M��\\�����&i�"v�K�̌g�`x6��l���*+2+ƾ�͘ʵ����l���^W[݈/#+z^��dN*�/�1.�M����?(����l��DD�i9��I��j~r��.D���!n�#�N>�����P�o�nTC�n��1�k���WPU�OI�z��x�F����U/�c��/��	<ÍT��ւN`��{���2�=_�������^���<(G缈s\.wN�zw����L/5�i��5:����V/dΙ(�ƈXo?�1q�o�=;�����6��=���j��������r[',���-�c��'w��9��_05
m4�'�D�է��6��6v�U:�!���K��Пջ
*[��q,�3��0��*D�q~����V�QU`� ��\z5sD�0i���t�ș��������M��uj<d�Z�d���]rL>>�:j���0��(V�/,��ܥJ�yc#BM*�MA�#'��+�;0�6���[��l$`u1Jdz��2���d'��T����3��~�3�9Ӻ�޲M{��;y������:�C��%����6y0US�H}P��9S����m�����������L��c�贛���n�r��~�j���u7d_(�Τuq8R�c�[J7�#����+0���S�K�ĒtG��@7��K;k��Θ�Kjxc2�sQ�^=^3��q �4���e�-�>����/{�<��H��<�؊��q<Czg�H��9�2?��m�E#�R)�V=qN����T�4#���|�m�M���2�׳f��u�Xr�ַ�F��Q�Ƥٺ%�?^N���[�鄓�^��"�w��^���{R��P�mi?b���"f��+W,TR�M�-Iyko��#8�q�ܓ�{X,�g2�cE�O��ԥ�����hl�,$���*8l�[����~�B+��h�����ᖖh�#�Ass��Åjd9Z���\�VyTN����Ok$�ǎ�?��hd@��6�c%��%�K��cKS4g��M���_��x�AM�������y%%U
o��~yw����'בy���p�jF�����-b����毗=1��%ԟ��4�k����sJg�X��i������ͷ��@\���e�����Eh{(��/�X�9%�#a�a��i5Aɗ{.�M[���U����4���gB�O>[	�t���\�
�4��r ԑb}ހd��o�2����g�Ś�u1��ؗ��$B̜WI��.��
�u�2�<��E�tw�������XonX���Pe��a?vB��k��2����\��ꡃѪ]���<-�6]�8e߿�-ʺ	6&N�[��q
ۃS�b 鋅~K��bޢ�=�> �ݵ�Z���~JD�KjjAG��{��6�|�d�i�*p{���g��
h�E�_�a頬�/�2�(vl��������߾��X�:�W�r���ү�^k)���H(��bu��k��5je�Z�\e�zsX�,e�O�nѣz�}dݼ����4�1|��t�ǩ��~B�&u|���/��_��J��,��~W�6�՘�M	*TP�W��Hw~��%T�FDw�#gt�� =F�כ*�>��2�l�_o�F� ���~��ʏX���w�I�����SA�
���u\�����}��hB���˶�sh/�	������kF,CpT���9���xB��� e��X-��r3�go*z�nN�Kq�)�ѧ�}� �?Oܳ�Nu�`d����u��J?��!�eaz=VnPQ0(������i7?@�!���%noJ�܌��e�yk(:��`\���9�d���r��-�����i�.eޘ���	THS��qx�kX�����2�im$�LƦLý!��ݙ
hm4�G�r�X�>��TJ�k�.�l^���D������Q�2W����nN1�wj��ё�]�>2-^1|�l��W���$Z��6RP�8戮��Y�
��2���Zǉ_�I��8�b�s�|�yj�~.�	<wH�SڱϞxd_�9we�A�9@�9�$찑�ʤ ~uA�:��V�����.[��Ꞔ������Q�4u���gXt��`�uE�|�v�sy�>��l��NNaBT9훾Xf]j�h���dߛ�J�%W�LoYq�QL��6����M��V��7��O/܇�R�9�6�B��#�)`ErL~B�ґ^8rێ:�̿e�5���Gͤ��u�h�*.�6
y�V_t�P�TG��Y73w�����hM5���2|H��$�Q��W 56���t��ڀ�jȔ�,RY�J_q�����1�즿�����l�ighZ��H139�`�����ԈVQ'SYq�h��5Nn����k���e��Aj��ҳ���)�����p���[Z_��p:��Sų�a?�w�@!xѯ�~x@�xA'vw[��f}�Z�W��6�2��=��5*����TIpn/��_8I���ZI��LiPJ[y-�����x��|W��\���\�H|�KD�9��yc�+g�t�� J��Zv�V؆qW��y����-�{N��5���B����N�{Y����a��>��=�����l�^�R�� WS�����Z��a'�"Y�U�����Un"G����5V(\��0*"��{h���[�^�ֳ`ꜫ��'S�/PCy)<W�9�O��
��p���!z �8<�A.�q%>�D	2U�H�{_/ �������1��uU|7�H���W������][CD��������_X�~ӽ(���VL���hڹo;��t��%bs��ْɚ/��{�8��?�y�׷��2=�`��r����, ���M�'R姹�;����O*�2�K�5�����T����bSM����o#��[5����3qɌΉ��j�-�-�9��ֹ9P�Ef�BMҧ5�����hfJ�?&�p��ï0j@_�&�=�˺z�\	�U�����i�b���)=͍��<�a����ӆ�&fyw��<�������:�j[�8��%
�W�aJi�}�]W"S�/�#I{�1�w
���H��i�#X�36(Q��5�g��;��MS��S�.��[�i��^�17>�*�W�q�pz��'���2����O�J��򴴟��9���߯��W��1Rp�_~�e��Y�/����b�/UUq�<V[r��~�J�]|�A�7�����r��s��x��w W2v�N�OZ�������"H�#c��9^����'ph{��`�u�2pk��s����v��*[L�|h����C?��S�.��
���Jf�L����L�w����1��_�\e�t���Y�XU&�pkA�O��;))8��)(i�LBg>ǟ��*v(CE�Ӈ�P%��i�F��⁁�v0Bvyy��� V(/"@���v6����q��;"3�J椗�F>,�M�SغQ�c��3�dӈ��a��9��x�}!�0�镣��C�"9%/L�n@�+�!Z�s�È�Ǿĭ4n�}R�c���Q��ĥ���ޗp�R���Αډ��J����X�P�N
��B������m��<�>��:ZZDttt2}ԟ��nz�2��Ne�|��'Wn$�%�勑%'ߋȫvg��,c�'�!�n:�,^���X����r�)�I(,q����b꩏ÞT���������[_)"�":ucߣP��E����B�دǐ�6G��ˇ��N-�l�*�I�E8;;OJ�S��8����������y�?�����)�Y02�P�]�
�����u���1B^��m��}��k�NWz.E�:j�~m��@^>+s[uS�oii���D�z��p�̈V��r��VY������w6��i-:F.�"���@ծ04��!�@e�W��%������*��6��M����3�?���~�z��rC�|�<zws˖.���N�]�}$���X�sCt@�n�@�y��� �����ku���_��]q@�E����!Q��6�k��s¤|�B�*y����~^�R�'�/OmΘK���
u��*�z�I��J��r���F#���>K�|8�b�/�����f�����C>~�dSW�8�ع���N������5�9�:j�_L�l6��RB����k,������[�x͚ۏ��`��9\'ؿ�jT@���ԴM�D�rʄ����^��mM�\�VL�w˖:�59s�'�C,���U\��7�?������ZX��\(��{b�DYT	�^�6��5�=���Xu,���%�ԉ�2)(������ɥ��*�i\4df���'��<<�(4$y,E	O��Ж�@�7A����z>���M��ү�*ӷ�aG31o��z����� �u>P�gh�0A)?�P��<:�'.���'��˻_�vf�� MG?`r�%�ٲ�ܔ�ebL���I�rJz����!�g�_$}M�s$� S�:�u>3��ψ	���<�qo���+�5m��4�{c$,��861��|���)򠸵�g���p����C���Tܾ"��1Q�J��B݋���R�+��װ��C<?�_C� 3���%���է�:�v��I��ݻ��0&���R)_����@�I~3�pN�r��2�n��Q����VR�#B,2�������WZ:M`���g�+j�NtT���p�3??����ۿ�Y�Ͳ�S������(�Rso�h�2��}��x���\��B�%���~�o8ѿ�s�F�o�o0p�8��DP�K�;'ocJ��lҶD�p#à1ݱ����s����5��\tt0a2�hȄ�8��y���eT2�,����A�P.�C8�I&J����j9:j�{�@g[8�����Wg�a��֛@-"gg��.�T��H��a��s�h����,+�,w=i��>��v����� �`�w��{aCn�|�>��!X$��j�R�^_�e~inn>�f?�0�=�Z1���$�[ɸh[6
��jP��@�����S4��):^,��5������T�[�(8f�:&�4:o��ɜ�G�������8��l���������\�j������󆝰�A�L�?U'bu�!�>��H���)-�7J^mo�S�0�n;��8����F������׏�������3���S@�����HS����b���2�r'�V���69�����ʯ����խ��4��,�lI��0�q;����e��,#��v��z�ؚ���U=���VH�1��>�JBӨ�E9"�1���O�1uj��ɛ�^��ĉn:� `v�|di���(|�������'_�o͔� �T�|e�@{�LY)oI=����B͹NN�u���ޒ�������4��w<���������������2�@�I�+!T�������C�w���=���ze�h2#�X��,�F�݅�-���Q�.��D��H�ׯ7��m���7�/��eS�L�,����]��/(��� �|�|�E���+�w�J��������v������P�<���_�]�~�/��s��5��x�7m:i�P�P��\Z~s`�#`��F�N6��c9<�nn0�%�ܑ?�{ak��Q{��_�*:�9���m�X4$e̚�H5��fHf��g�ΘŲ`�U�-�.`�!�v�ɓ�Ց=�����������޵���AB��E������������_�ޟll���)jhh,,����bL�b�X�:����8�u���@�^�e>�-sj_�g�.��cR��:���Z_?��,i|Y:{��?�������6��6~�`P�7W'j��hGZ��
�����;ao����B�_bW�����������v+���������k�p�,fo&��aї9�����%. ?����c[�-m��Fc�;��_�[މ��X;�R�����"�R�~���K���������}mov��v`s�@�J��9��oo��.����9��ʜ�>�"u�B���+�J6!u�+�w+����W�Sȷp>�<�JP��x
[��;�jK���Z���2(���}�$V��S���)��f~��^�n����ɸ���3�=��bQ�^��>�qb�� �bjF۫P D�k�6��kZ�<
ٕ.D�5cvC=�����d�/"�}Y�����[Qɔ8͆88�r�XI���U|&�2�1,�RP�����
�>��i>�#E.��؀���z�ʧM�U�~.��K;)RJ���1����b�ڏ,���qνec\�c���n���P3&�1�Ҝ���\�2�j�%pJb_�u�{M@�ʔ*�������4Y=�<�?��4���y	b��5�������H�<�p�|H�s�|��v��D�wvt��� �j�ϴ�f�� ?�_ҲI`��U,q����﬌R�UN����?�o�s�|"T�C�i�\Y�w	��V�81�n&Bٔ2��5�6��	R��9��Ÿ@����`��G��5��ŵ1`#�d��h�K{Z�fA����V�Dr`ܙ��c�T����OJc����a4�Xm�fƽ�r9��y�*>́+����g�&�g�uǳ���#+i&&YǃqcUs�@��S�\�"U�s���7���&[r�o���@� � p�2�/�ӛZ��������h��/�"��վ�M�ٍ�@�r0y|D�۽r[2Lv-rQP��#G.YQ�������ߺ� "�s���o5c6��~�"A�O��Ȧ�qQ�������tqU�_SJg���PsF]C��I>�k=�2L�D��0��K�'�b+3׃�\�nT������P��-n�7�b����E"[�(2�Rc�K/w�?K���c8L��@�����}4�8�e����3Hz}�+�֭!�� ��Ds�����©;z;��SĠ(f�`�]+WlƎ��H��G0�
T;Rm�hr� �g薉d����0����K0�蘧�$J�:�@4o�bnC��?K0U�FoV���M��@����~�9#M�?��̄Eβ����'|l��M����	w�9����{� ̰���OJN�����$1]�THg�)U
�?7�6p;W6�F����`�+b�g�r�ǭ-aeUȏ����KWg�!Xh*�fy+�&���|���{3ڹ�zΥ�*B6����4*ս���k��'����	�˅��/�BeN�fҿ�ɣ�3�4H�D�Y�| u����$M� �������wk��]����$G`g�����0�(F��Px��p���@n�>TaÖ3�P/��ɡ�d�^���6�����_ƕ�_y���G�3��� r�C��,|ϛ��w	��b8YI�Z
$"Q��'^7�X�s��Cy�	.�,��)ۭ�m�Y�$ޤ���'�(��]v��=��\��?�x�h���b�osSKwR�[z��$�������������Q]��sZ�^�E&�<��=c3E���ʟ�&��~��o+�ZZ�39�[�6r
�tDD�>���oֵvE:�y+bf5����}^}�a������/7g9�ƕA��n|O�|90����r3ʈ"��ϝ�CP�՘��q�3��w�y�F�՗�x9M?��v�6H�O��N���Z^�Ϙ0��*+%�Z�`*��K���P<�C�:�7.�;��lĤ�Y�Om��1�O���ED0�N{=�m,��u��k�7�ρ;��__���
p�#!�t�����Q#�2㖘�C��"{����_���JO�u{�9x�ɤ�a�����W ��5����Cp�Cp������ݗ���K�]���	�o7��^=��������眾�}�)���<-V���C�p�R�0��`3����g@��g�,"��/�H8�����$�J������(���He�Y�nv�"\�8e��,{e�5d{����7�I���
4�n��@�����Z���w�sҺ���_�؄���I�һa��I���5�l@:������?�6����I6�߄O�����.R���7��fbS~-�f`C���do����k%t�DR�0y�f�r���@\H}�N�KB|�rv`n3N.)��gf�q�˰S"�;��?�.Z���#��r?gB��:�.��_���w~�*!Ŗ+^r���l4B�{��0�Q�Bݞ�Ľ��m����gƯ��b��w�|̇3W�Rm�9n�lW>�F�!*�w�&~��}�ڨX����f� ���h�q��?T`�LOǇ�e<[����o7�LW.�����������nñ�*lL�Ӳ�˽��Ł�/	�p6��p`��z&�7����y��k	�E� �A�<�FƟ$�Hї ��(��+��B��B{�!�ş�33A�ӵN/���)���%Z9 � �5���iݘ����R��kU��I!��Uӳ 27-Y�����5��KO���ޚ��\�UV���׋�#�3����J<��3w��Y�+2p�#��%Pr�5�چ!��vKO|�8��֧�6l�;�ZlF�Tr���fI�	[�B&g��!^FW{��d��罐R\s@噬C��뗆Dga�:I)�,j��)	��;'������rw~��+d��g:�(�1�����7l�|?���jo����cc�ǹ/�J����r=�w5�%�N�DW�nȺ�������PY�7(7SGkʡ�l�c���K	a;�!�`S1hw��m�*c�0ºI�J:\i�u$g�x�E�Z� �r2�#^]HwUgQ|:���!e�Z�p�3��q`Rc
�3pV���)^X�рb����f��?f
z���ڎ�5��w��*����8q��u���m��Ib$�niiD; p�]՗���|t� Ff[-ߖ�lX��4����?���CY['���>:��ӵa�@Q�_.�35y���B���g�L�(log���oJ��{�w̨w�$*��ʐ�n�PW4)IV�f�V����_'w[�����m,��V�>�p�l����D���J:R���W���7�B<$v�/b;�>���~���Х}��W���o#���5j�/��N��Q�2\�`Zx�����r �'Ț��AN)4> S۰����YfYa��MRc��t�ZbTV�S�}�h}�a(�e�~ȡ���)����ř?�CU��!a�8��H�,�]��2�֨�����qa�9���K2�D�m�:�t/R3ݛe����"��:m`����
��_-�g���Y$�����Α��bv��R7;>uc��� �7@����U\k�>��ў8���Z�;ߴIh�r�%���A������-?L���;j,/,�V�E�'��ӕܨ2=~��h'+��g�Nl�?l��>�7�ܱ��W�P�DCC��;B�<��r�����4��hDJ���>1_~�5hM�]k`-H�m�΁�	��VS��cI(���	�� ��I�f��W^���)��G�_J���g�ڽy|������� t�z"I���{�����p�����I��t%D+���ҡ����O�}�7�o8���A#iK�6�C���*�\��&���吖����Ď$�����OeC�O���|au��sc�\)�a,OGL����m4_W	9�,�ޥQ����Bj�r}��e�"Q��;(��o-���|+��Z�c�����%��O��YX�Z|?97X�t�a�}�>1u���R�xk~�4�ޔ��)t`�Y}JCy���X4#�k���i��_�Y��0R��e�״�4��Z�!J$/���6�L+��n�:�o6 VB��!�(J�P�Ł��)ѿ�:��ąg�`���Q�"�0��G+Ni�h�zl�S�!�%Ov���5,��ŊC��P*��uo��]�<���!�Ǘ8�V�����6#��]]K����c ���Ku�^�'��ٙ�n������^�R�ꏇ���3�%��E�tv�B�Yr>��Q�Br��
x�`��9ܪd=��JTdHj�/��c�������v��t�P��ׁ�u�۱���!o��eN��--5��V�[zMw��QS����K�w,���I�O�IO��_�W1XN�K��t�^�U�Ώֽ���*�]������L����b#c�����v�fyb��ٟ�2�:�4���f����X�=Z�������@
�,������(#�]��c�^`�zR��`����7���QL8�U\PŷN��!n���O*��Y�>�}H��z�I*��=< �����-?k��$��x�/����]���O���s6�J���L?E���8��
���? ����wƺ�cO�5��gLNB0��,(���	�ׯJ9H'�i�w��0�#�>.�#�%Hn�n����|Oօ����#��啿�/�����~�k�X�>����z�����h�<:r5��ǩ����~�h���+N��+��ǘ�!�qcI�:܉䤏�a�4	����V�4c���C�;�G����y�!���X��y��{g��<���|k�U����A���,����ȞVD��s#��A~�,������>�j/�\��Y���2��OtG�ዧ&�>Gse�{Y�NGe?��e���@	�����Uu���i�LF��v�9.�B +sVY�lR䉅N9����h�!�G?�7H�P�=L8:Y>�^-�ZW�,v��е�8S�I����깛��[�����'Bt���Fi4��כ�U92���f���Rdu�7@!Ô\ta�?�q��G��w8��<9I8ć�ꑰ�l?:IB
�=��΂QX��0�����N)t�����j����27R�-͛0�I�c��;�M����,���s�#y#�R�.�C��&��r����&������c�?]����mѽ&twE)Z�"�(�g�9mCT4P`^��h�5�/����ZM�Z��-��E?'Ӥ�^��%��dt�M��N(�|i�q&=�i�$V�fd8����_��:]�ȉ�},!��hf0Q�	�|/��S�w�ǡ%m� �@	���qxtr�ޝs�J �+Bvu�rc�*����q��[c���6$��EMY���@0�����0����/w[j�y!j�|d�r�2∌�Ƅ��F"K�DQ��_��+S����V�pF\A`��	���D���ջI�T������<`s�ͷ3�B$��w�:*#��O[҉/>�ŪYf)`֏�j�\�T~�1QQ�G�����f��o/�W��+
�p>��[��m�<k����x�L� ���)��␠�^e��C�V�u?��\�k�D��t�pe+�\�����*y0�W�c��3�������"���i�d�R�~�������+�1!ŗ�grY�K�:�BU�Q�Ws��2��G4c�N~S�L5��[��($���+��N��Q��R���m ��x��f/s�;�O\<���h���n����#��� ?���eտ�`�JPs��ԗ�tp~X?�ܰ��,c0��K0��!�� zˀK]��+JĎW�|�b�ss�2o 2ڧ/C^�](.]��Ѭ޹ɢ��ӂW���u�0=��l[��Og��wv^�8���`�Qv�؟���\`��UCzP�Ҍ��r���r�#�k��H3���9����2E��'~k�@W%�SLS�}ZᦑV"`��6ZS�u!��ߠ��*�f=�������~'�
�A�@)�k�F�}��k�{���؋f�}�H^~v��U$�ѺN��D#[A5��5�Q3��C��q��wgt�v��o9u��>��=-E�/Hg9�u���.�bش�fE.�K�!��ŀ|8-b�7�X�9�j}�˖�������"���*�EG�؅�������2L���ˆ���߆"U?�%�����ᬥ4�Q��/��rPR�qq1-�W��I�y��TxY�p�����6⚧#���l�k?��T|�nk����P`�]D�2u{���Y8D�d+a�i&k���F3D��T��'����	��.w���FB0gJ���j�
��2��.��*E��G�\��(o4�*U�z^o�>�Q�����
����O��K��6}�ڳ��9�Dl� �2��󅩹U���0½�4�Vces�5NgY����T�Z�ttML51%\�Q�nRe�KXbᛤD��x�s��'��q7G�,���t��3�ճ� ɋ�=��PB̩Z��Ω]��=՝|��ԭ��T�������Iq���!4ԙ��2d�0c�-'H�w_�M��Kc�wsh��cZA�E3(
�J�)�0J�h}����5�`#8ӑ�M��"�^�|����t�x�ǋ}��b��Qk_?������055�}��}���=��^)��y~�1�jYQ��U�P�r{����KKu:]%>���n"S��ݤ�HN�-|����1ٟB�����ܵ	��gXHG���i�|�<4
�~��u��iA�o׿�2�#���ޞDy)��t���Y��!���62D��?l��o��)�� �Ռl�ܔ�Z9!s �qZY܉�V�|��eL�u���EIw�v���姵�m���� �F�-���X`�ky��+��]UK�_��/} ����o��/��8�gEo�'�vP8��sGt�!�?�I٭^�?>!w�co�ih\v�.������9�����$��#��f�Њ�0 ��%�1'a+�*��]��"��W
����IyM]�I	9���c^�y����EE�J���������33"������~��@R,�,�۝��`��U�jD懗�h֘��9�v(�Ҽ}#?
Ӽ��#�7Uţۥq���z1�5��ֶ|��o@�	���X�ZZF���I�Y�Ʈa3ӈ�غ��o�#� �����J���n|K�O���?m/�X�����y�|��s?�x���;�aҌ8��d�S�ݭ>��Jt���,F8%p�
��=ɟK�aխ�Z����jT��`�n��r�pn��/�κG�΋���qޅ�г���3eBV,��ֻ� ѺWɝ������0c���3�����ď3|���鯛�v�W���Ъ���GCN<X���k��{q�##�4;������}�e9@T-SGI��;��?�V�Q�|���|��og�G �Q����ew���~�=/���X�hx�o�O�lT��N��ۅB��`fј�0��Pղ�Y�=�Z����^9C��t�LߙZA+
k+Ԥ��`�yY�B��[��-.<+`��D>l�e��N�<Rl7ٴ$7�<[�"�O���t�Djc)`$/�'���4I!�%,>~]�Ce;���6�QU���(X��(7��T�\!N`�U_~Q��������3c��W9��!��6���*fI�4�7�>��n��X�����>.�:|��)��������.��W���.n�w�z�|\���`�i
�|ҫ�dA�����0t	^$���_N��l�d����@^ir<�װS�E�(��4�4��9�w����s�_��:(��b"
b6/�_uUF�^\z�珮���[���A��]b	gH�.4}po��ܪ���n�}�k��m������0�5�����s"�:=�N1�6,�Ҿ�`�v�g4�y��yl�N����_!�,�s
���3͖��S�	X�۳�����5�����ι�uo��[���ƥ�՜[�Nn2��.����EV��_��C9�Ɨ��H�D�Z�LL�'o�d��nd��O�_p�w��bS�r��}R�4�7FE�e�{��Sb��ik��6�\k�.��*oC�������
�&�g��������.���N"6�G߃��jy��qk
-��fw�?(��P�� 0(�u5�k��iw�,��D�꯰Q��5<e��I,�Y��6��<z�@�A�LUM-��j{�đņ��൘e�Q^�</��\2�a-E�a_
u�&��0�B_ߏ�@x	*���3ysSy,	#RM����/�`���BKl��+\�t��
��{1�&5[$�z��ye�l�:]���2�vp$�Q�O��0�}��'��б���6Gǽ���~���ʇ����qM�o>P��F-!p�Y�W�H��`�n��'����ΐ�1���6����A0�~�H�I!N�uҨ����
�YQ�򡘜V++���UV�k��շ
�&+����� ��$�[������&��(X���U���Eu��B�IL�O�d���j�PC\XQ�j�I9|��&�l�*L��Z���n��ZN�j������
�rՖ+iH���w�6Y�a��ly�ȹr��A�8*����]���E��h:��K�H$����u��Ch���(-�]��R������D�N:��*QN��s)Rݻ���%�l(x�ߟ)��wvB��A?c�2d�do��u�::��qs�0����Ǭ�~����&�Ƅ�3�n���[0�^�:�_�IN�X/aw���y�#���Wn����f�S.�Jެ�'5�������\f���wG�'��y��q�X��oOM���Q�����,�����N=pE�Br�~�n
]b>b8�i����s~糷G�'o��b��o���^��Ja�&Y�=�k]^̾�{�@�("'��˭z"ڭ��ߚH�Ρ��ɥ�sQV�i�����q'��}�$��[���ף���TD���c�z���}p7�Y4 {BԜ��o�v��~���g�����VJ��W%��jߠg\e�Mx��)�����"�RA��< m���@J�f�A��h ��W�ZXV��(�"|F��F��B�H�9r-AD��
꓁A� �����R�>�vb ��b�(j-=����޴���}yFp��N��d��s��M[%v�ַ72DjPbON��)k�DT����,E�H��=�8^�t���?�R��� eQ.��/�eN��N"f�����2��+���E1��#���'�H轤ω,�*uJ��Y�*b��p��vu�3���Y��Gfꉽw���n�0�[#�8'vs�����}�ý�H�` ��m
l�:�S�W�.o�	ѷg"c^��4�H�D�T�d��ѕ��$��ͷ$��H;�A��������M8�4zH�K��g�m��1 _�u�{�)y$ǜP��q(k�5����l#�V����y����H�́1����V�����@��@�|�&��m�w� �����6�;��m2[0���B�5@nln&~�Ɣt!=:�-�`M�H5��16���ףF�2����]#�hƑ�iu����588���XJ�WN�w�gνʉe{���E���@ �9
�&�\MC	����PCn��r��J�j�B��j���zL�����[�(Ur���)3Wp��R���u;>Q&c(U�(�w�.F"(�{
��.SSTt�9��������^�e��P�O��Ӹs������ޞI<��#B���QZH*�j����$�
8�,öe#L�R�9�%KKP��	|?rJ̈� '�ٮxgN~��p�]�X|O\e�ǹ�p}�j�W�}���:T�QZ�%��uQ�}�(��!-Qq{/����eMǰ&�z�-]�e������8�X�ˌ�|��`�<��(�jf���^$i��#!�����Ʀ7��^�ˮ)���e�:��bBPwwt�	��7�Qv����*0��"0n�&#(L����N1]CbL����bTV�}�f�I0�}�R�0�3܊�P~�EG%��R�:x$UT�G+��ܞ�ɪ%�l�i'X���U+�,�21�Ƒw�ߖ�T�X��L��3��%I���aq�"Վ��UR������͐>:��:�t1��~���k<l�&��.h.0h��,i~��#��N�4�Ir�ΖZy�671J��A6j����H���n�4���և��}���Yjp0t�^:�i�K��&��L㧬��i���Ox̪Rh�Q �.�.|6(> W�p��hG���=C��#����@mx�5'I��>ё���9�a����ݟz���q����Y@$��p����چԣ$5��1�z�z�}#n>��i�@UC&W�RQJ`� ��#�E8�����&!���	��������	�.Q�qr
�z�{�������L7�}�?�ǂ�@@�9X
�����s�h��JgՏV��X�����M�'�#�'�9{��ju֚C�!I,,[�{s2P������Ć�U�X�̉��+���
���Oϕ/wRP�����Q�_��*8S�BS�U��b���P86��� w���$��'Ȍ{�c7����⪨XQHu��7�o����C,������J8�ǔ��?���VG5ے����0�LM���}D�?#R[k�A�'�-ނ��E�����G��72ӥQ�̇�?���Jl
cj�i�ƨ��m=����8�q��@'�[���~v��	6��n����C��p���$�ؔ��|���ӣ�����] -��ڊĞ;ؖ��l���.�HtCҸ<R�4Wa=4@*_P��Fm�Q��v&��SK�I$�zg�P^�n"����m��r <�h�"v���/�`KwBũ�ՌTfw-��wҊ)�~�߼��W+���$�+cq��ޑ|������;~����g�{��}]3۬�#h�'��w��s{���)�����8 #�R�
�t�WW��vQ9�x�¤)`��$v�mL8�{g�$![��{� X墲)�QTS�9�~��צ�`����T�lgDϏ���AF�0��
ط���k��c6�{���`�����������/���.|9J�4�r���Fb�I�Me�%:���0����r#�])��������F�{V�����âGӭ�5�V��;hk9Y��hnۦ��E��!�g�,��>�o�2��Fʯ�G�>k�:�t��Nnմ�L�[P�]��3ɸ���a�p��߮Tօ�$�q� ճh?��+i8ڟ(����$PL��G�_{�^�i2~���(��G��Hw1��S��ف�M��6�G$T����b��#$ 0�n>�+͒Z�c�:aݺߚZ�+�{�(D�u��|U��YF$HO��TEQGR�.kE*�+n�f
ڟ�t�;]��h���,ڡG!�3�\�.����dn���;�<�֫	�:�'��}q��߼<a	�Ka AQq}5|�&ܰ)M��H��DݻS[A� �:���Y塕&�/���̀�o�������?�Z#�W�ۍ���|�����eO���?�$r�M:m���"R[;I���0Y�\�B'��$9Am"Q�m�'h",fԥLA�:��D�δ
e�/��� ٌ���.g;�T�q%W�OU'�O}�8��.�c�yn�����/�13y6B��CU�Xi5��#m ^�@� ��㶄����O(����J|�iWL�c�ۦ������������p����w��Nz���1�K�����E=��}jJ�ǳI+�f�P=F��ix{j�n��
��*��~V�KFІ���Z��뿺�c 7����^"(y�0�r}g�UGz`�����Nvu%�x.��a�����p{���6�>8:2>�~����8n԰��ķ�����g�5��! p���������v��Sk�z�/_AӦ�(znQ�� ��t,؄Mx�ݧV]��p��K����p�_��qҍUT�7��Fj��0XF7 lߓo]��r(�3Y_ޝ¹�n�l�(�o��چ��]�@�2Z���({rf`�2ع�[^|�'����O�וE�a7�c�K��k���@NzX�6Y��9_Z��!ߛ�:�ڙ��W�hy�$Í�y<�5������Q,������k�H��}I����DD��b������k�u�'_%$�S��P-!�G�] �WJ��~I�c�/���1=T�C���8�J�s�dℭԞҠ�v,W��<����Ϫ��e�����w���:��ᄢM�˗����s�rKI��C��Q����'	C�C�s[Z��AUϡp�Sx�S��Vh���!�.�:΃��:���-�8+�o����#�Je|�P���dl��ZH��m��� 3/�0�����m͏��y`�G�`�iz�!�KA����P�����<��"qC
��q�تP�6�'�8O.6+�t����]S��UI��XX�Γ�ڛLd.,'
j�j���E�R�t|���xN��kB7Fq������MQJ���dI�Cgc����~��k����o[5���AA��sZ�u��)���O�9�$J��P���A;��1��Tp��B&���0ݳݤ4��"�k��2�+(�&�2��Pc=�����A�	�wn������F�U��O���.YƳi��#�r(��/j�o/��r�6Y}6�Iμ�	�n����a�U�Sл��B��╨�&:�`�	 ��<kF�?ooo� (��d�J�<�lo`B�6���󆤽����g��"4<>ٰ���7���B�ͯ�v_�[-�F�|��u11s�Y�6N���B_�ⲇ������Kl&v��ˏO��F�/+0#����a�/��M��]�.6πgK1�`f�+������t��0f?�)��W���Ĝ��~+T���}k�ة��8�jB�`��2���9�N�Є<d��z�s��}�Q~+:u�5J�d���5�����-��r/�ۅJ1�\�[��0�*{>�_�M�������5�=|�i����~1���af�Br�(kX��̍��E��oѦO 8��Å���P�����Bm��(�������X�1�����������b�Ht��9�iE�\���:|�T6L-7R��_��^�,ry ��*��Y�����b���u�Щ4`n+���6j|�t5�ͦ>�6;���bz����������{m��Q&��H�z�7
8��bed������u��ԁ��l¥Kܥ^Tҷ�5�����(���	bB%�$�
�,j�3�z%v��Ln��:@���??�б��ڡ
�yP��)�ev{REG�T��a�]l`�`4�7�PzƋ�#��ԏ:�~h���df��w��~��S=	x��#�g�"ؘȖuH(#�c�P�q/�����@��3�	�c3� �q���gX|���%�6kZ�����Q��0������&	�����<dt�}t���y}�~ˆe�uy�Y�C�8]
�SΤ���_R���w8v�?!�(^�]Z5S�8V$�������[��q����!�@��Awjv9�(񕏦>R\r�P%��\�[8�mA��I*��У��K�A^_��+3�^����W���|쭟-��&x����z>��)�ŀ2�@���v!0 N����5�������C�[��J�Ou�:�o���H5���X8�Y2�'��]�L��~�{����j�Q�T)	�7����:�jXQe�K���YF�����m�+�kV�z~���tQ"2o��?�M5w��Z�.���~̞�{�H����ݎ^p�	�͇�>�$z߃���f�̓������<�@)s�/ vv�����B��8V]7������Vԯ<��D%�CA���%���X1�9�c(�՘����e�o��eLI�AnV �oʫ;4�G�.�?�Mn;�9�*�R��#�=何=<#�"�?>qpSȰ˫�j��(� &lr橡v#^�RW�]�����b�����Vح�Q��� 9d�A�����R���)6`m����Z��%kب��,
T	š��LT�(�KaCp�|�Ҵw�)t��;1�J:U�8�0<�S�R_��J�aD��o���q���:��U���)��#�4�Л#�E����E�x.��,%8u�S��7K��|�N�6fS��u\}�Ex��K�2h�ҳ��<܍%�=v�p���lli<W��u�p�
[h�"���+-a�;[%�������G�:�8
�~�n2R݋���T�Aq6�=���ȃ�?�I�|��믏�	�Y�:��%��!�fk����c�?�֐&�cf�-�5�-U%��1�d�iF�����fW�k��(�������\Y<���N(/g�[������'��W��; ����ּX����v��W��o%���<�yo��]g�V����R�Po��att��M;8 ��qEW��>h؆���r�����2m3w���C�zg9k�$U��.��6�R�f�`���~1c�E9ǌ��F��V��qKt�#j��iK�N&��Al�h��(��,��Bʝ'��^@��#�B�&&�o�?��W��jQ;D-]���8 ��N�iZԢ�w���Q�`�Fq�^Ծ����]<��3�S�����r
l�(����4f�i)��&+w���@��
2&5 m����)Rp�k+Lc|��(q�O���-B0�$����F��D�p��~^E	������x��|z��(�$db����r�F��AL�Zh������`E�v�`��.l�=*�ָ�ᐠcg�c�4��z�E4#/y�[��e��1�0cӲ}oH
�'g������N$a�p7Ζc.!�P0y��D:nѷ�SI�*j��-�G���n���|SbZ�iV�8a��P����9�CS��*rH]�~N'�>e��Nc���)�$� �`A��05��w��3�*+a�@�+̣e9�Tޓ����ͷ��8|Z�pc� ���6~�W�(�0����U碩Gg��[�875�G�c���d�8�d4��{�>���܀N�\z��a%dd�Z���~���U��$���M�_@�u�~9So]oS��7�xXS�9�8�+��~���&���zp�w����Q�TK�����Y"HN����jI=��0�e�$�P�5��U�⽙�d숾R3`'�.k��~ �����d�b�����隍-���)	{R1S��D�x��^�%&�vf3���QBN�mHD��f�HB�߲�f����b�~�1^ �abbG��@x��l��r8xAB'
k+�?{�jR��<4�R�]�zR�i������0r��F�r�ǡL�f2h.�c�A�e{HF���o�F�ϥ�=7�q�g`���H#X�hG~��0D0qC(�f_x���Cu�H����-��*D�w�D`�ٰ&���,$�@d)�7m�j�5�l�kE�4f?������Jx���{?��Sw�y{����G��s/:��2�FDA�
U�9O�}�ĩQed�~"60n���IB��cq�'o��i	SR�S���'C~������/��� '"��� O��}�CIP�Ƃg}������p�5�=ݝ:���ה��%$�H	H�=��>+�����鉌<�i���A'8�0xi��A*TT��H�g�gl��i٩������D����}�ȯ2�o��{A��+Z$0K��� <�N`����;�hӷ�K�i�Q%�)�X�v?�O�D����6�k�	�����#��w��js�
�����ӆ���a��;#=��8u�r�Ʀ��7���ɸ��5	�%�X)�	ײ��`Z��;q�RI@j�.Z����,�����y��t��}E�����|"�u(��39�>.�����&��0�X~�IX��:^����\E���E���_nnn�
rK��h��Y7�&�3f�c�����DLcV.��!�`�h6�>��h�4����?���\���v�����Y�.(hv��3	Y�0�)M,g��L�_�Z3��B��8��Uܷ<�3�+(�3^^��������:�}%�~#�n� �K|�a�gэ�@I:�T��vgSֳ���t�D����w=J���R�'X\1v��l����_�u�Ng��Cʮ�̏��}z��;(���o���7�vҶZ�� ��9���h�S�z���/p���	�gfʯvZ �f
��뻦&������=�ôQ�·��-킟y�	-N���'��}�1_����z�/��}�_�'�w0�Z��b86GGF������0��n�d���4�?��4k����k=�;XY���������8bm��0l":�ݭ���X�)�ל��-��22];�z7Fw3I�������PͬϨ
����B��G�Ui�ǩ��Y��	��F�%�K��0>�M�Z�`/�?ru���y�����Z�z����N?�f�.r��܅!J�-�5�{�Xx�[��,�G36"�|��	~~�/��6��_�xx?��W##��sarS�������$D�����2�-�]6k"P(#�f�m��[�����0�=0��{���$����R�t��&&�>���։�H ���bu���i{?ʫ�Ӥ����l�3:ZI9鵠;�z�C4����~���Qs��.�&���@��Q�l�H.�yHC��%��& D/���	��P�?���:9 ����\Y�+˜6}oɡ�j�hZ@5	���m����J�# �{��?��wJ��%2,��#(��"\.��?�>��!��]�Gт2�f
M4���%q�H£�1qˤv�U,�&d�oiP�B���Z�Y���㛀�� �����>���tY��Of��q���>55���b�� 0�P|Yh|>�@?��\�j#R�_�L�7k��W>�J�8޴R+�w����+�{xNi�xB�JaL/>|�Io5��H2vz)U����MO�P�/6�7?g�Z��� �p��p�j���)V!	Rd fFp��?����w�����2v9�mD��D`EgǚP�^|�`''�+�\�N�x�٤���~H��n�C�*���q|_sy����VFFO���v������ب%.�rFLө莽]P`z��+��M:�Ɋ�˱�P���٬������]m����6���YN,nU*X�x�ؽ��]+�(�C΀���/��~��̂�k�ݣ1���cvn��!�FQ�e���`P]��C����5A�䈓�OӦ��(���(֧VcJ�>�
��nm�esA�Q�͍rt�ŵ��	�{ew�ljW�s�<��E�G��O������EyF27���j�v�b����
���	�EL���z^_��0vG3�������~�)Dk�T*�i1FF|�K����`�01��3�Z-��4�$4�3��x���W,�l�� �V����a�g�'g;RhE�5V���뫒 y�&������*���J�g��W�y=*����X(��Oo��G���X{a!J�ƹ�F������-0�Pnl�]p�9G�r�qc���&Q�[�������p�/vHG��@ο:��zN;`s\�R$��`f&(������U��	G�|������A�����sk�dH�T�Yѳ��h����l�B'R��͖�im`2��`_\'��ʊ1��˭䀱�fŠY�>l�����ߔ���F�����(�˔1������S�#H��ͤ*T�Ȼ ����d�j~N�����S ZkX�!?'t� �[U14Lh�]413�������7z��B�X�;����X?7�����&��z��Bm.2�Wr�[�.ΒV���zz��>�@W*�G��w��g"6M�r�a�i� �e�����7e��L�Bn��D���ʩֱ|��P��:q%���щ�N1�T���q���E�)~9/��o5�pm�p�Ϟ@�%���"N�+��8�a_��^���~u���Ѻ�S.kE�x��経� �h��Q�[W���U��ce$���m#*}��ߗ����`�-��%�"m��[s=���!<�b�[�OY9�E�R�!� ,s��  bH܀��!2�1��g�������jx��a��5r�1D_5��S���j��ìL\\܍x���m������әx�7��>_����][54����gE�o�7I�5�ꉢ�Z� /k
�a=Ůڰ$?J�{�(]��&� Hz���t�Ő��*ä�KC?�'B�����(b�DjL��'��!"iS��Ϥ�'*��3�2��X�U�@�Pbc�%t�u�)�Kw#�`N���IM�ZX]���˫|y�8��9[Qx�Ho�<\���P�sڐ�1C���������f���Q��Kp��� =�/r�v�A��,�Sڑ�!w�������|Y3v�f[ږ
��rX�\�h-�S8ևs�rD:9 ;����([]����hl3��̡�����nM�p�x�zo�v>����j#�R�W]�)m9��Db��	�sN��蕚��Q<�0.&6�GN�Ȳ�Ϥ�����Y*�
fh��DkcK�y	GG6�]�999�2�1X����G�~��L��+��Zt�������щ ���I.GGG� �f�7bC�t���*D�xޤ��L���/*���dѴ���<=���BCa"8|�ӂJ��YHt����5��x���O�e>w����lcp����)b�Fp�DKf�~D|db�4P�쓍�?7��4A���P�B&�~�#a�^�q�,@��䢊�f8 \`nn���ڽ��@ӎ�U;Y�E��6׫�b���h��%�hj��Gg0��__�X9-�Z�����kT8=_����I<�j��n[�a�����>E����lQ2��h���lV��H�=���Ÿ�]	\F�p0���G��=\;�Tت^T Y����r���ݯ���&�1@�K�����}���#��]�6��&|3�]4��2q�l�k`�FE���s�yH�&\��,��:�hli�l���m��!�-���ڮa��-!��Hw�� ��t#���ҍ�]��i��Mw~��z��C��Pֹ��sE���5�F�33��R�^�&�!�ٜ���o]��*B����I���V�B�u)��d^A%z���f���Jk�D��ν�SY��B�Td�r k��쎑Q�bx*��2��`��Z��v��8��_��BY�Թ���Z�p�2_K�=���{����G���d�o+��\����a*HK��zg˾VYLѴ�nD��3�
���'��=9����oo�oDJ��y�ϳ��}Lҳ���s�YAMB��[W���4l��ݶ�(�0?����W��%f�W �"''��X�����`<4d�勥ا�Թ@��Wʋ�s�����	ּmq��Q���*�G���ŶE9�[�{0�V���_�E!�y�YD�R�A���*�J;��m��rm^)5���H��ތXd*���]}Z�ԑ�9�/}ߗ��a==33���p��Mt6�Xaަ��6��?3�U6� ����$�-Sհ�*��KE����'撴�#N!Kb�gL��j����M���0�đ�m�ȋ��Ig���#W�@��nP�'��A��q�ۙSd�;݀Á5y�X��R�f����~���|I����=��$C���_9qJ����hMԼ���d�Ywi���84$�x��'6��I~{��"M���)��d3RR�ْF���%�����Ȗr���@���a�g�?�LP^|�%����K2�����K*#ww���Q���xm���U��p��p$;��Sp�z?|c�K�|_�^�d}}Q�Y��F��2���nw���R�Pa���a�/�K"ڽ'�]�5[_����>���uCT%[F�F�ݿ���f���3�i�|���F�����&?ur(HduY���2-��X&���(,����'�C'���Hl���O��W��I�-���(E=<��AUm\BWxF+,5\��b�
�[��)�FL����uk�͇�����9Q�2������5�s5��5�:5&��'�ĒVlT9��l�/p6\0��ب�Ă���(j-�1�-��c`��Ы��y�V��;&O`���[Q�r6��M�NQh�������*���@]����j�)�J�J\�����fx�_-(�Ωm���:p��[��Nn֮��e�^ł��;�}E���]�ll5�pr�`Mm�Q�Ɲ4K����vO�Q��a��=����Op��}tq�\��%R�?4-�2��f�7�*�����b[!zhhG%�7\�8�62ߓ���L����q��:OA�����ֱ֮2�v��훹�P��(��r`�}	5�7���<I��BC�l���9�Ρ
�e��zS�E{H�\^K�Ͳ+٣��!3��aһ{Y �s��QQW���mK���9*֨���)Tb��0�{���!NsɆG�T�?��Y���$êx�-N�
��À�NHKcH�j+VN?R=�o���B�Z���ұ�鸿�\~6{#vP�o��4B�#~�+ڽ�/�ʔ�T�?-��*#����{��?b/����+%����Mvӌc`Sly�Dh���xr~>��p�gY4VvX�l������A����D��"�O����������s����
CKY�|":4�N)k5���aq�ט�v�0�R���i�_�p��z{(����°������T*��h�C���:�ۿ-Ҹ�9�x]�ǂ�1�,��_�w�{�:(�Jٯ���W1�TC��AE�܉��l��!VA���0��yo�����SR<k�����P}��d�o/!��u�H +=��r�5�Hݤj���V�|c�j��dD=Z��{��^�����K��G���S�~f馾,#LG��G�|CCJZ�1�"]�G����h=�W�����(����?�����Wl�����Y��q��8����%���$4u&��eml�>��^z��G��|��$W},���:}���ձ�9�zODA���>R��'��x��&�a�� y�0���-��}W�+�p��x��Y
�Yq�ڙ�	k��8�2{s�'�T�P;/�����ϖ<����7bF���5�Ι�fPU�wQ�g-��0���1$�u�gR(�-v���F���{sYD��U��6�hʓ�Uu9!��6lE�䲚 7�H�O�2�����[x�k�jDP����'f�������r�
�mw`�y5C�:�9�R��'K����L���
c=�\��R�O��n��N���^�&z�����7J�t�Г`�A�"�dq)|�o�Y�\M��Yt	XM�A����1ٜi��Q'otDvw�P��ʈ_Ζu#�y�.l�A���?t��!-�	d����"����KP*����w)�㜬��0�����``@�Z���5��_҅���S��Ư��ğ�\LX��H����+HR�b��
	�yA=V�XAH��pz���'������h���2�C �������L[���$*�Ac��B�Tє��J����ug4�l�(v}���y�D����1�T{����{�)��W+�����(����v�o�9j�ϖ;�����ch�`T\���.����Q�y��e~$'eP�Z���瞺�����w�bY�Q:S���
\�v%�T�sRW��g�^��GO�
 �3��Ⱦ�/��^��{dU4�#���g�z�ՈL|"qB[�7�^u�'17x�ј�dC�(]���c�cX���Th�R^���nF�v�rN)��6�q�����͝���Y�$|ߒ*o�`L����>���
X�~����j�5�	u��i�N���HY]p8�I9��?.��®�AA����k��H�P1��
��Ȁ���m˛����o��!�����h��)��tI�Ĳ"��E�6x����W��0�����G��EF����Ʌ�����s��%RQ�)!vW�&���:��-R��I�K*\�)��b�leM���sz�B�f(��,/�ײ� &�z���]��b����n؁/�l����մ|0��ڴϚ;�j�C��:����:���|�
#5�nh�������gZ�E��bU��$,��%�q4�+��F�/^�Ew ��|�B��4���uW��(�ę�ۧ��u���F�3dK|���oc7�/[$]�w���Fg�w!�v(D/�'�o�嵇��(۪+	[��$-CD�W��4]X>Y�h"v*♓;|uV�<�%��-�,�W�iJvv�5�)*��V��7�Q��'"� e) ӱn���tt���t(��ө� rc�Yϥ�����1�D7�ĉz k��v0�w{89�d������2����	+�$%�co��w1��WW,|=�����#�a�kL	
�Z�͉��@�._"xd{e�y��G߾)2�|��􇨼��Ak�c�gA~Hg0�nXs3?PjGBBB��%ةz������p�f�K������a������E>�z���\���Ѥ3�������G�)���3{nͥk��Hz{��TipDD���èV�o�l�x�`�&�M:�e�F6�u����)��Ed7��0����\#9E�X̔L�Gm�)Z]�N��3n=<*���m�1^|�U>�I��f�G�0��V�����~�}gTI6ߩ���}��ۚ��\61��<�=|=�H�0r�I��p5�2�6#FD�k���R�'͍ĵ��ROBBH������g��P��T��{?������%�GW��G�@�%/����8~�'�'ˣ0^��C����~����D���*��I��1q2��(ގ`�:��r���|i�LD��쫃���n͉V=GA>ը]~T�p�͖�dȸ47�E���� ��2�2�!8����!q������Kt�J�Ԁ�mKo�Y�*��|�O+E�`9W��yҊ@o����\䊍	���?2TeO�ДU��b��I�<���Qu�r�`
�]w��i�$��g���F|���ϔ��>E���WF���	��~�DQΤWXlPN�5
Y�A`�N�������Sa�� d��!��kj|�=n��ӻ1�|>l*�t;��H�9�1�pg#�4�r��'���ZHb�ecTmЭ�-�����M�,Z��ap\E���>�$K�~+Y��ѫ��'>(�񉶥�������I��r��L�.���$m��+��{��cΠ��ǝ6�J�����}��F�������v�N#�wz��/*%"���Y��1XIOOҬK�X��`�C�ݧ2�i4���:!���[n����h�	�؃ϒW�N��r�M�B�0ޣ�]%չ��p�`�|����8q<c�/[�P�_��ưP��~��7�u�A�#���q߃&ei�^�%?�@i��FN���������F8-�!uXS��<o_�#�>�]�cQ�E�r��������aHL�~���>_�
<������ W/��pԨ�h˴y� i�lon������꾫�Vv%�IҸR9i>�bF��G,�eפ����XE�S�������MJM[��6��%�����ֵ�X���>&sO���������3wJ������Z
����K����O��0�/TG��	Жؕ�R�D!�1+?M� M�QP}-�����,{���;<�f6�1�|Ԣ�2��C5���s���ۓ��÷�K�Bi�(*wͼ>2�_�����&8p�ս���ۨ��r��~�) svv�Ȫv뱔S㨫��΅6~�=l1�C��2��cͩ��`�vr����4��I[�Nx%���=@m�df�T�nhP��u�]��g�@z9ɵC�Rbe\��w�>�ٶ�?C)�m>X:H<�o�5c��ÌW�����ۂ��c�7���F����Gd	{�:� ��qy`x\�Ƈ�����yf�l��}s�x�{�lڥ}�}�}su�Q��KE��;�����+��������Du���f4�B�ѣ)��_M:ϩSK�2��F6s����p�dd۠Ў!��v���o�7~�H@��Gr�^�O/k��W�%L�~s��ߞ���WE�;��}_��ƴ �[W����+0�:K%4B�X6^�f�{�����#Ô	6nV%�W|}@�o�;Ψe��/#/�a���l�VE5����\���j�i��3OG�;���\6��S���j.2��u�_�/�����w��@�i�n�*Wc;��S�B��[E�X�����vwBlvw)��#&�Q�%��l���{��3{~��;�vE��۟УRNm��l��t���τ�~6,�~]c�{yA�5���؝�3���}3�՝���>����d��|�G�-
�! ��']sܪ�&��@!Ш*+��V�8����e��7vk�A�+$��F��&�H��<�mݠ�hE�W'��P	�n��ݻ˔�}UX�"�t����8�E�-���B5�M����O���g�@O_N�(P6��C�CyʥDX�y�^���
���v��!"u ����9��MOOM߷7�/7?P��G27f�F �p��Up@�sj��b���FB�h��.kEhܹ���dx;�t7<�4�����w6˞��Q��{.��Ĉ19����|\�:��E&��DL����>�=�S�p9�X3�+���8�1�ڍ���<ߞ�	~C��+D��֗�pz�$���x����ߎz�[��ټ�A:k�� pg{#��(o��6�E�CPUd��,�i`�u
zS*W��4v��_���˂���MT�&gf�ّ��X�9�3j�d�>�ܝ��l����%��	�Gy���x�6xG���혁O�q�u�ȫ[84�	�rrJ:q��Q��x@f��d�����	�$Wn����%ڎ)����S�^'�n��L��-+���:�)3�idE�!)˺n}Xn�4cM��4��di���)�	����.��� �-�ק��lv���^)�ڰ�_��$ �/�)]ۚ���VP ՐׅT�}���n0~ty5?�a�F�vye)��A&�o����N0Eq?�omoǡ| q�M��jXv!�fi�Aɟ��/��z7��&�~p����V5L���-�Fa}	�o���bɋ��18��S'�P�������k�׬��d`��*��I,�u$��<έ�]����e+��J���7�3k��J<��%r��X���p����$�e�⽢Z�6!ɉn9쬶��4]P�b�������7�h\V��q|��·=�D������x��y�ײ���;J@%�С�᭠�,ٸ���ڄN�c����9���țm�/��������N�i&w�i���`���gՖ�y��@��ƛ��á��?8��(�o5V�\5ҩI;%#㳇!��3���GF���}L<�a�q�G!��pE�'������,�D�%�I�z3Zw�hE���X�c#������0���l���#�D�:��BK3L|��!�DR��*|i*����71|��� i�VZ?�'S�Ղ�/V���� t��Y��E�ƚ��#���j$��$�V��2G��~�(g�����-�hU���Ig��������إ�C���_�)6G������o���+�-��p0��xYUx	�x�����XZk�U4@i�ڙvd�6z1�4Q�Y�����#ƐI�~���)9����o!ʭ���.)K�#4��%�_��
�w�H�/�P�,��@n�*���9������,�q������4\ ���S�©����k<x9+IˀґC���3jk���� ����pr�7��g��y�a���ݥ�o�g0�q Gd���u[Kl��*��8�,�q蔑�Q�T��ˍ\"��I;$�H���s���-A����@Ә�!��j�&��5`E���E�D�����_�)%ipp�F�!"0}"E|�3. �V����rp~_3p�C��TE%26e;[��7K����y�ڛw7IocW������C ��~v��J#V���_�W������YBV6~r�k������+����(�&K$#��-R��jNY[�pb)�r(� *�e���C^�zݲB��.�O��-T�::$ ��:������>�3�eYx�6xW��eV�������^�M:��MD��1Mp��e�7�;o/�@S�na74v%D��9����D��x*�P�L�S���l���S�~u3^M�1��Q���Կ)Q���v������sO��-��w��
�t�U[}�5�������:�kX�z#���s�{�&yj$����4b��b��ܴz�%��4�K�B�@�-Eķ���Zr�@KQ���҆��RD����N� U�y�e����z��]������}q�K=�DZ.?/9�VV�z��X&�~9�vۋ����@���0����-��^ �D��P������ɷ@O::Y��~b� �Έ<���oH�\M��HYk�� E�>w�z�"w�·k���LG.�LDL�Z>飦Me����,��|�~�!�5�a��2�- ^�o�ݿ)������������L�t�p-]�m�v��!�Bs*~x���O�PQl��CG�J(Mm�&�\��\�[���`}īt{C��	�;&�0R|�bWO����c0�htwk�PZ�T�\��P�P4��L���ח{q��'��z�њD�{��9hEXI���d��a�ex;��WM�5�`�̖�6�t�_so�j�[����H`T����ͺX�F����k)w�e>����tpѤ΄�(O�����+��]��ȴS�s$v��{�^�q+��uw�x�F�M:2R�"���S���k9x���Ǡ�z�c���%���5E�s�M����}D�n34������`$^U�4��1�(�P_��k�M/��b���!-���w'Xˢ���1�3Y�aĨf�<�p�d���c2Ǝ���"�e�`F�eI�i;��~��h7s$~��ar����e	2��I �55��v�^ <:5�:K�갔-��'AC��--r��D���
 51$� � �{�F˝��ů���s�z���t)Vn]\�����}fk��o��/pm3��VV�i܊��t;3\r��JP�W��u�dϧ���@C�԰�5r9�QNi��Z}r�k�r2��9����[���i�ZH���Ϻ�9~�n�c���c3	azϓ��B�-3og�������+�j�����>�}��g3�(�n�KoC=���ݴ�kn�a�z���V��%�w���5��|;�&����僋�$c��z�!��e�TOc�����7���G.�_Omu~���mm���B����"\�����T����-�WF`5ޤ��Q�=.���D2�~C{c�.�;���:��b�PJ�iE�g�C.�.��;�J�K<�|A��Sf|�To ��!9
r���S�A/��tI<&s�V���&���ӱ��B6]���="�g�J��<�@�iL6�iy`��M��
~m�"<,�V��f��Ygm ������M�����z`&g:
��$�����?�C����rc��ܓl���y��y�V�4�C��x^��m�|��h��1�sR���*!Uo��I5�kj" ����W_zy�	�
���v7�b�>�=�/�Du���+����T���ۿ���Ҭ��)���]����,���i�[)�_dQ�+� Z�T��ifό���ܖ�XE�����T��k,�c�ǿ�������?,k���F��C��_�5 K*���4�ˌ�RG�3.b�H2�S& X������o��
G���`a�*����0@��x˿���!�����������-�2���?�M�7S,Ny���#��춏�R��r<O���ߕ䬚���p���n�g�PR�j?"�d��v�z����HcŽ�QAR�[<�}x[�|��: Q��ܻ��x[9�Y
p%e��(�%�l�8.�G�9�0b���MQ�N�r�o�>{��D�JmLczY1��'�> ��+�7:�>��4�v˰�B���x��N7X:�I(�q���`�K�\0֏�I'�绺bخ�#���?���%n+vǏ4a�.��fS��U���?�mT�iE�$a�8�47�������N����F��;����ᴯL����Y2���߸#`��
�w_p�>>�?+���x1!��������u�l�n�3!�"46#�x*jWFW�~����X�Ku��k�1��qͿ�k��LhQ��nN6ޡ����z����a��k����P�Yo�$�I�ysZ8>8	;��o���e�ܤ�ږs�)�s�W)M�`3n��^!��	�Zi��sc���3�av}�r�k*��+H�wk[,�b[?x�6��p6�*��
E/4�����:D#�A�K������q��[-��P�n�����"P��G�����,��(Dͫ��Ȟ�i_��R�W�i֦�2���E�XD}Ʋ~��D�F6�\h���2�n<f�ޞ�9MSɪ[idj�yE�+1�N����!I��>�x��G�e��*�;���k����gQii�(�j4~�|��Ag_Q�?[.fs���a��ĳ&28�U�f�ኛOK�5?��Io�vv��R�E��o^�h)��/��d�{�k冚>�U�����63@#�1�}>J�4�/?�WS���ͮ]+�/��\���x{t�S�s�$�yB��s��"ݯau�s@��l�W6NN��n��m�⾛_�«r1H*QLp0��ba��;�z�?-�o���ƯO�f���-���?���ډ�5�hoy�9%����V{w�#"O۫�q��A*2($�c�1I�rWv�w�x�������{3V$��k�H_���_�T��?z��=ݘ�I�@2
��;�����>���&�LSSfo��i���Jo1j�#����P��S�Y�w*�����|x�'�h�+�/�+�R��~�[f_�;-��-Ҏ���������ƕ2I]��~~#m�i��v�nk%�د�m�����e����g ���fY��d�Ļپ>2����r��5K�����[.������~�%	#
)zZ�fZ{5�b�T^��V֖b��pH ���oȼ��D�X�oF�T��jxЉ!p2�^��k9ra3E���^�4Y�~2��`��{p���إ%mm�e���?��	�f������#h��f��g�~d5�Ȗ�LϏ�r՗L�����)2�N�)��񜭞�E`aD����m~�c�;�z�?�v��jf�ǝԩP�G��cW}��JƬs���dt��7*�7��`���w�J\���x�)���~N��ӓ�����M箉������˩E���GZ�>FFT �6Z�ݮ��_y�GGz�2I��f���!��� %w�b�Q�P��7pU����d��&Q�&n���`2��O@f��p�e����DC��D�5���OD�g�1�����+��SV�GG��.����8�A,��	�ۋ��[��zӫ#�:NF�RQGGGe8����:n������}�ߜ��?����e�����H���mhÜ@�[�N�_�n%�ޝ?X��NtS��D*�ȸ��o T\����� �o�Ji;�R'VUS3u��l��Wb?
b�OJ3��&~���z�L%���/f'-�0�_F��!_^7n��!�t����R.?�/�$y�fȹ=�~]�.M��U�G�SD!�أ��M;v%?��*��J �Q�QS� ��5\d��H$��]�}�:�%�?�y��-�<@x��s���c�؁��B��3j͏m���\���Z	ږʟ���l⵬k��H|�L�%�c��x�5A��}h�������ʉ:]�J��s
z�p�D~<ͺ��e��M[��:��BEaC_��Q@���P)�&���w��y���%��1��DKS��,E(��h�&���_X�{:�-y�!A����tkcD��b*��"plL~��c��Z�7�.+0���.���Bb<�Wyu��7�A�qAI?���_?���|�c$H�h�x�]��~���l�xX�Q�����B��~��Y�,� V��6�#͏^Sc��%���/�ZC���J˅��j���=��TE�(ޑ"-��z*H��,b�����y���Mz�����e�b6.H�ңdcL�^HKj²F�L�5��ƃ�]/��[M���o�O⪿7�K��9���f�X|������t)Ywi�^"}S��,��"d�uq���t��a!�Ґ�b�\i��&�M�?i��B�ܼ�m	z�Y��ۼe����!�:4�ϴ���^�d+wji�Hf����.���x:�.�tE|���-9����l^������{�v����� �����?5H~~z�^�+���?��k/��`��y��vC<�s������C�6KWVQi�1������G���J�&��h�L:ބK����-�-��I�zL�w2=��D7�/��� mtnW3��P�P3�	���7hhhvw����:ff� Uv�LP��"�25bb�q*jQˀ��V�jОF�k=���4w��~a�~���;$��+�W�aN�\�)��Ĝ|~�&�m��7Vz=���I���K;v�W�o��
7qi��Ŀ�{�͙qE��>/D���af�j�l��Z.��_����T^Pm��37`�P{C��}�������FI%T�L�m�����l�䵶v���Ա��Bc�hĎ�~`����*��@L����6�QQ��!��3H��\���5��S�P�԰l�spx��v�� ��Ll�X"���p�Im�&��������8e�	7t����v�ł�e�:�"��@������́� ���P�.��!�*�q�`yc/�Γߩ� z��A���K�B��t]��7/O���n��O��2�)�%uL��V���.R:���F"ΐ̿���|'KqS9C_�H��6Oϑz����C�J�㢉���:�o�[=������\N����a���n��k�%ԊB�r��ףݐ���o�f�v`]�$�u��Y��$�F���I� �#��H���XG��<�)5��y�@�v?�mҹ��D
�N����3���B�*�����dϧ�-�-�1ҧ3�z��9~VV��mQTU5.��q�R3Z�ˢ��UK�Q9qqT���Γ�y��V�>�k�-3k�[��1�;��n��f�g=/p��[�^m��TM
��,YO�����0k-�uE{�Q'+���@F1���ɬ]�'s�����Q(�F��`�^},���f,�V�Y�z���&ƳŌRm3�Ums��Q��,;�bn����m+N
X�f8O���8ӌ�ͳ�!Ɗ�/�:�W�ג�w��<��P�jߖ+\ﵟX��U�l%�J��n �������7���G�[��~T�\(�&�N>�u��\��S��^�Iq�£4�_#6Ȉk�W� �=ڌ��ǒ��ya�h��>��B9"��J�PL��<�	 ��2[o���^M���GCn�ċ_5
	�ksRg~U-K��_\�W	�dȶX $�y\�&h����N���Y ��n�v;o�%ux\[G ��I�瓤��N,Z�m�� A��|{_��jC��ZG�^T
���D��e.�`q%��
���h'Tk�_�"?�0�rդ�=Bd��9�m�1|}�'9jU*d����8@.��qW����?�B�kGN���u1���Px�?ؔ��0YI�{)koan^`���o�e�3ۡwW��-�~��߀� ��AG&����V`��I�.8If@��I��<���s(�◣��X��]��a�����7���P�w?~�XK�j��t�����Ω�n��93W��6ǾQ�.�۵W	���.��-V�K�-9�00����"��s��x�C���]2>�[��ͼ��)I����Q#��-A�^]������
��J�Y��ۼ�Y1�٠x_��X�,BrUDU���!�p���k���i%�H$,��=��,n'	1+�������PQCp��I]]���W3@� a��>���0n�D��ʉ,1���-��qCj�wu�^X��5�^����,��~C.��7��ú�o�A`9�g����1�}�F�%���ˏ�tZv{�$�TUy��g��?Е��7�	��E���gy�v��'�տ7��_q�AI�G11��>�͙c5�4�5������)�u��l,�"�D������b�{	�]v����Y�;�y&��{d����^�	��{��j6��*��.'9kxɊ��
8Zơ��h�`S{�m{�;
�E;��Xx�4�F���>G�Ӣh��{?p������n�^�G׾�W̯�/���p�ll��Y��'�:� ���gT���,��e+iW����f�w43��|b8�^'��N|��9!X(����Ծ[��Ӎ��܏T�yC��Z}�`���R�Gw��x�q&'YD*9�d�̥����opc�{�����ٝA��ʭs�.z��Y�r�<U�\�럇�xxF��g��n���k���o'�L�b���`��y�Z#�P���E;R��Z����aP�c�W�B��Ph}�m��>�ڝ{�!��Ɔ����6������	�޽�򪫕onli|w�⏫~g�1�3,�#FW�L�{r��tnuAr�lXʏ�M���u#���3F��~f����f��`���7��K���;�ߚ]���C����O+�z������� �8u�xc���Uc��R	�l���hW]���l��;��j_�I;<��a���I�`ʠ-�y����pں�%�q��ļ}��{�g�:;����9熪�Կ|1�A�&8_k�@�Bh\��P�V�:��{Mۯt2�iU��v�w���,��(��\Ri+��~v	�SG4�J��-`R��	�����]ն旝r��;Ocj�2W�ObG�z�Z�lh��.ɯ�P@2���׿学ԧ$M�����ۺ#s����C�F��I���NZ��6(h���6x���s�i]X��~�2Z�`U�+�,0y��5��m�l�|<�6���"N)U��H�?4����șc��u�������R�l���]�ź��ރ��б|���7��:vk��m��0�T�Q��y���&C���� (:���-K�j%�PW(�v���ۣ�jܝ�o�;�.�>	��L(�4z�x�[#�J&4�G�����ɜ��}���Pu���\��M�.�����e\K��
�Kxy��8�Ɉ]�!��q��RB�#��x�]�������s]A��'m@��`�� ����p���̿�ڭ}������(�(gk^PSg��7]~������5^e��h�(�.���JY�ݹY�zo��	q���y�s��-D� 2�R4�!K܄jz�|B�W����W>222vP"��r1ֽ�}u8��Y��Aj�������% 7�51���*毴�׶�U*�+�-_#B�eׯ#l4V4�4�_Q�s?ּ����j��g��s-����Y��=�p n�3� ��Y�I�Vz�%�Z�������^���|#A<ߩ)l�>�s��g)j�P�ܰ�����&��4?��?�r�/#S��>[�����
���5I�Z���t��������;�<r��w��#@yꎳ��w�I�K�}�T��k��>w�m7��'}�:� ���hXhYk1�כ-st�V�ش�K�XJ��ҭH��S�u��E�ZL-ϐ�=�5E�q�$�#��Kc�["|�Y�p��F+u���)���)�q]��w�x�̧J,��,>s[q�*�z�m����yI�j���r���s4詄��p�� 6*iߋ��V\R.�����0aj�	䥠�#S�Ma�(Ĥ�'���0u�h�i�i����u`1�5�ԍ9�s�.���v�C�t��v���g��t}Dd]?�T�w��]��{��@u����ZJ��}ȶ�<�Y/S��0���@[�!2�˧�7�<=��"���1�P,�%f�rHL�.���'囗�>���q��u�O$RPV��c�T����t/eQ��"�Ъ�Ҕ��ɂ�_	ǩz��1+w��,(R��L�G��,�Q��7�2���)�Mv��� ��!�'����w��O�Џ#�b�(t�r_<~��s���3Z�j���z�M�8�ֲ����.?
>�nSԫ�ok�ds	I�{���s�8���WM}���q�L�r��*�G�ƀ�"N�w����WN�M�F�JP5V��V�̃s�v�^^$�aʒ�˓�p��@�0�QL/�,�������ː�h"�[Zm��hN�ۭ7
w�{���i���թ��	�O�!�_2Վ�y����B^Z����[LٯI���W�(�]?J�ɕ�^g�v�EG�v��i>sC��[�R�Wr0Vs�ʞQD�*a�0�ı.f�a�UB����\�A(B�m�вݠ��b��|h��q��s	]QJ��HΩ�e�t���t!<�����f���`CO!��,9���oH��>�-;�[��
�eEٚ��3��5�ب��Tux��k����?`"�ݨe�.����Mb1�L#j"B��7�+?�����q2���My�w� 0����/<�4;u��>;�d�a߬x���Q>���걞fY���������J�)#ݣ�A�x�'��0�a�t�V���G����'n�����w�x�q
�ە��d#O������ߝ�m��<�"�8/�_�@��u�x��],D�����coF�=�����Le�"+^�?oD���m}C�z�W�1�K���!�@Ϻ+6l+����P(���I`?���K�ͬ��u���,q����1o��]��' ����@��3��%�U~!��B����\{`0
BW8��[o8���QmQww����a|�;PfZ�W��8�@A1������h $<���DC��<+2}���kh�N�<5����4
��d�P���H�T�]�Zq����C k�J�� ����f9��z���w�JU�t��-�~ �ӕ		�z�5(&�K�[����BP޴C�#9�L2�z�xx��BQ�{�Hg�X��� ޢ��8O��7V�d/����:���Q`g�`^�����=��A#�T��0���mՃ�!]�'b'}���U]�fީIO�s���Q�KRc����s2�U�Aʯ��}�'"��<���"#���z_o��WEb��C3�pť��M���J,)��P��XK;��Sl3f�6�J�PH+p�<�cp����{�Y�7$�u4@=ojյ��h�҂�N9!�k����ݡqzӕ�T�]�-��3��튲�T�3-j�����a�,�K�������t������KG6���X�� k���p�b6ƀ�sR�ˬ���z�V]��K��6#��ф���x�M�Y�����
�3m������Y��=�TH]���y�څ�d�2=�4�ғ��6�fD�~hWⓉ+�%�(k'�4^m�%M��D6�\a���0��	d�N�J��k͑$g�X5
�ݞ=���-�T>t��ǩ�����4��_-@�ɇ��
�Ƌ<��6� �n����G��G�B�PP���W�ܞw[�S<����q<+<5FX�H�����E|w���9��ef��!>������-Zޗǋ��n���GZ�5_�� �Ʀy��:�!�����C>�X^	�;Zx�%u	pB@��D�yi6�X.ő� 1�s�Pr~������0�?�v��-�p�c?��=����^4"#�`�0�<ã+�:����k��_���])�qb�5�O�䕆��0����hj�{iT
�{�n�1�o�;��G~�`���C���p�~����P-v|��jQ�҃�DM���@�=�1F�~�q����fw�Zw�i�[z��5)]�7��y��3N��)��E���#ꭣ����q@:�� "�ҍ�tJ��tץ�A�����N�KHww�����~�\ֺ뜽��<�̳g>��!zz8.RZFw
ؚ���=l�S�=~�ؤ���ViU�o�(��[����Z�g���65���ھ�?c����֨i�$;���K�����WDxڷ�]`�<W!i��[��o�o��9S�q;�P�0)�Wz�#��j�#���YA��$a��0b���M�{E"6���&K��Y��t/��1W�tɗ�FbU%�����)�C�,u`���
=>������o�)F��cKz�ڰ�ȶ��d�	�g \��� _�]�n��X:��J�����_�)+tc����S�ɪ����Ah�x���dg���]`��R�1�� �B�G�F�������T��0�w/U��g�|p���,
��b������`� 益��\��7S5TK��QȂ$�>����D�Z�ϻ�Q�a	>�ɳ���E�i�}��'����%fWa��,{����`w�(kDv���	�K7�Ph���޽���A�^�%��,3���6UA��Q����^p��ڞ����L�iJ�j���Ep�@~�A�%q�~�Ulls�7��u��t�T�(^���@x�Ӏ�3�:�nz��`�o�@���٩�����P�(�NM��3�\���L UpvfE�A�i�5����sVK�@��e����0��;�I���g���=We9�U ���8S�Y	��X�/5�'�V_q�p�v�L�|Z5:��s�¾;0��8x��~K�����y���Y�����]���V������?u�\����@���������6Q��w>R��\�x��\O��J�iڻz��k[���0����E��?E����W7�T�2K�F��cN"Y�C�%�\2�Y/�^����Q��UH��1s��i�?�~-z��E�{���w��*`�l�W�_����.7Kl��B��J=Ijj����|���Ǝ�ǖ�������ɘJ��@�U���N�p���d�ˉu
z-F)d�v�{��c���F?U"5�c�wZ��1~^nL��#B����(�V�T��:bOp�fdg�-�[� �0>Y��ip�l�������
���$���}P~M���*��d>��C� ��K9Vi$��\kS��6c��q�A{���&��ǜ��<�e6�މ�ы.�ĥwgV�t銲��GaFҭ��=$�i-	�+�+1��p��R�>ެ�oɟ:�8מ���F����l~t��?�}7I�����kv��p����x�4��a�|�c���{FOI��h�����%,��S�gKGr|�x�m�me���W����h��?=+��j�t�&�{f�}��B���0Qz���'*�EuI8i�f
C����0���%���j���L�>lĈ+��@�xS�'�
&|;���5Cy�9�+:>.�2z���w�=Na	�K��;PDv�9��_�E��z'������E�O!����.y)�`��B�~� R����E��ܠ���D�\�3�e��}a
l}�$��C��f �]�R����=�����ԯF0cv3R	�_&7u�]���Ven��Wp�찒�<�W��:stKR՜���C}Z��$��Wz����v?��E���_��?u�}�|9Ϛ�!��O�׶��Mnz=E�;u6���ֱ�;컨ٳB )3�S1���|�Z��ˣc8K�2i�e�k�o�&�'����ir��oS�}�lF���`�ɀ�a�2w�`�}�VR������jة�w�W�m.��a�>�o�R �;;>!�d��+Y�_$""�����F��_�P�x���P�L�-���kQQQ�k����c6²b���jf� �V�/��ퟛ}8z�j;OF��b�7�cX����������%�1���;���ВXO�A�1�mZ�������׼�1b�6�}�M�|��9��6�I��0`�>��W�BYNm�p���HE��l����i댒�Q�O��*"i�Ob��|��k�����������Pii��ь�
l��e|f��	�J�Ji
7"���|��(~(����UC����܈��������E�����e`��
��^Pцr��	�{�q| mp���m)����a>�U�t�~ӱ)�
|7VPLd���K�E�������CV�(.$w���>�U�@s��H)e���$�a*;$���N�	�%��^
�rh)Ƒ�g(�����@�����z��i?��ؘqѡ���1����֙3F_+�n�lti���]�=DCMm��I< v0}�R)�\{|���?5�4�C�qؒ.���'S<��ܘJ�N�]���cE���2F�]�s<���^W��H
FTL�\k�	���,�|��+��$� K���mi1B�ii~>�Pr�뺂�$pf��G6���A�iȬ�FJ
�T+��`�n��vzMU&")���/�\���L��#�Jd���o���<�ҷ;�!y�<D"ya�'��T�qC�&����C�bF3�����&+����S�G���~�!�/�h�H�,�$����Z��|�kz_����iX;��b��&�ƪ'E�=��x�4��eV	U.��mQ��̗�u3��K����=9m��ߔ1�Z�p
�4(��f�Y[s��`�X�h��-/\�Ea�jq�� ���4�]`�S�k�M�?f�Y#Ѵ���i<g=��%1z��|,>Vk��X�P�>�@��hAj� ���b�G�U�������ƒ�9��ׯW��.��γ�w�������Ҫ��hR���P�\BBB�����o��&&Vu����`X H���z[�]���^���}5j^��8����|��U����M�ý���8&���5�Cw�Y�8#F?7I�7.�1DXIQښn��Gy�4�]���~ge�S둌����(��"����U?��b�����9�4��&j!��nu�[V}4	�$J���_H�H́���es��8�l��<�17	TI���[[[�}PN�䢟A,�MU �K��$>��D�׳���)@��~��d��R��VY��*S��͠��2ER��Ҽ����9��\�D�u��n�̎�?A5�k+%+�/G_���K���a�/�L�c���⠳R���GU�;�ýB9I� HUW�����<'� @F�����*�������Px¥�ځ:�՗wW�<3�A'k�o3���c�̜���ol.pjFC�oC?GT�.��L��z���^�=86\�a�W�{uE&"n�X#�8��9�H߄q�5�=F��ڳ�~���]�a]�E���z����)$	��X���7P�����g6Rw(�x�\,�av���xR]�� �o��
D� ����+@�*�H�3�_��kp�˜x]�G��RӬQ��s�p�hr�{UC����AU��~��d�wKk�����m�K2��s;�o�>��|�#��6|�nUg�iv���@�'C�<���Gg���d��j�n���]M*��iϼ�apĮ��f��}�t�
Q�ZA%��b#������}��0��׹�kc��>�V]x����*�������ժ�m�ݖ^S[�K����丫� ڲ!k+8=|��*�Ę�:�9��3����H1e��$C��8�8�q��f����?��*F��پ/������ջ~��]C�����c��S}���2\Ҡ"�bSF3�5���DE���>�-��	;n4�ݭa�eV��^�n��5�V%D�9��� r�|�M��Zfw�Y�N��']�:)�+���y�Ar1���;I���E���9+ƛ��(�z�
����!a��e����n���=u���cg���jwd�ò�_�n7YЃms�{PG��G�qs��Gr�ˎW�<�ʏ�����£*�_r��Լ�ڻ���2 ��Q��Cp���!�&$H�g*���
9jW!���Լ�b��+Y�
zuU.F Lk:�<4���&����e�6��g�	�}^O�j��`*)Cc��.YQo�����2����}�OoKqh)�����۸n(�;�ջ@�~v�\gE6����Z�\��us� �����q|D[���?��Y��o��r��<ρ:��fqG����e,� �	LH�q�g��-B$����k�o�<J4:ƨ̡�nʴ5�b�!�m��ݝ,�}���e+ßBY�1�\T>)	�n�5bj�;!r�/-���t��:�^�|�����e
,g)k�{2ތ !q%�L`ECA�	y�#-�Ul��®M��̈E�V�x��
�{��u���\��jW�4ݤ4��l,>a	b�DP�j�?��v`��i�����a�^L%�;	b���Q�ӚX:��Z� �D��/�Ò�Ҷ��99��U�L���D�eK��g��܆�!��!Pk1�mX<���p7�k%jj\\0Ĳ��
�������������Y��*)Q�;�\�� ��旰�*�9�q� v}̢o��y�6l�Xv����jF������]g,��U~��V��bcq��9�iz��]�]�Tn��N�wȼ�
M�R�i�9V�s�dΦ�\/ߗ�u6��허���+��Vt� �,��%��вM�]⎻���G�[�ʹe�Iܖ`r�+�A�
?��'��[��y�<�]�B�[�ފmD�IX�-o�-����~�4���2fFO�3NOWf�5�lU/�N-*����?/�Ő��A,$H�Qp7��10���I�c�}�GQ=�Pʬ����][W�z��!��PM.������ʙXx������9ˌ���Ē�V�!妖h�nY;}��>:�â�;����d����fd���QӤgͳO��Y&GlY�-'�C��$���7�8\6�N��<WB���݀)���&&�`�l�.�D��Qf�Ƣ��OWB�d�o0*��3k�K��A:��`8Q��n��^ ǭ�� x���O%a+uZ[�*�z1.#�]{/"@�G�hĀog��n���G�OJ�������R�>F����A:_C���<o�"y��5D��5N��7M�0����c �po+��8d�����,e��X��A�yϩn�@"U��F�� ������:_���z�������<�De')����f�=�>֬�e��W�#��#i��.��Q�ߤ�Q�tϚ�l�O���T*̏L��\S�ԉ�~\�Fh;-	Iօ�c�qp��G<Ǩ����"�g��52�蝖nF��w.>�li��U�
��������9��wn�	zm\?��H������ߜ�`����O�m���|^3-��L��Fh����{��'�(6D�r��� T���s��4'��<{v��q��)�6_�e��<<_�pE�Z��7xm�z�[�m/Zq��\i�/�Z���:��ۚ���g߽�$f����F�4�1��Wթ�'��w�?��0���r�/�ǡ�b
/���ql����=�%X�ݐ����j ��|Ps�Je�#��;�Ɛ9�`2���R[�)�tm;Qo����~]�4�K�K��eA�E��F�-_���3�{ktؓ�����/W<���	g������an�De� a�n�fJ�v:����3�,�	�
��;�e�����~\p��K�a1�cyL1$& 7E��ވ��b�@/"��&Wg�D*�����t�k�}{E|]��*ŷ,r�l�\W�H��Yq��s����q#N<<<�s�~�7g[`9��tcp���B�b���氤�9ܖ/��	�TH���a+W��*��I,�a�Y���텣�KY�֣~��"���&�9��(h��#W�R�+�.��Q^c�b�H1�8��tAf2!%L���9���R���"�Y�;��+2�r�4Y<0�Wʜ�߷xP	�h����T8�����D��U���>�^��<�
>�� FTe9���*\����7	��%~���`�A��jwߨ皵gQ�tP����m��fq�,�Z��xA5X��UX���[���+�����c��>�90R�,��,�D<��u9&���ѣ!ٜ�H{Y���A�����>yzt����p��^� �c�J��� W���+�?���Y�1}���s��Ou*�����CG�y��y(\����[q����
���⦛�,��)�Ex�����I�F����x�q+Nu*L�jX	��4.��ٱ�Q��U`k_~��{��u �J�,,]��p ������ϯ|q����>�y)�k�����m�s�"ˤ}M�"�,&�;�
��,%($��y��g��,�?[NMz��3OM�8kE*�a�NI�Q'I��8�P���אE��
�&�tm��(L�
&Bg쯹�V���		6z�#��T���ޯ�")�_p����	%Ѩ��u��N�����|8��h�ݛ+��*aN�j�/wB���5Н"�r��ؤA*�O$��)�`����(` ���
*@6���}ç��y3ב�}��%is2���Y���s�����5m��9��F ���᲻�u�xj���o�EHct0���!�
�U�ڌ�
e�NL�P�r���D��=J,Q1ҳ�2P3���XA� �/�03��֗�E��!$e�9��[?w�p�0w�
 �z(Id3�� �uX_������w���3�M�nG*�d
{�Lu%ŷ�%ă�|��!��:-&�R6�/������5����LÍDF$�߬�d��k��N8���\a2��HW�m��H1��㕮_Q��j|{)��KPC�f��k6�Z'k�`�7Z�Æ-��P,�݂���#�t��$!��G˔ �_�[qo<���I�_�΀�h����;fl��Qi�&F`�PW_�ih֘�+��]����Aٽ��2ϒ#�$�F�P4�w�g\�R7�z�K[�)�8����Fv�"6Y�o&W�s-Q�l$�
��-����>o�GT��ſ���趤��L����u�N�%�S�u�~��]���N��L �V?[��:��R��s�$R����'�2�y���)�d2Э��#�'����`�N����E�*x� J����6�aར�U�s$���|8a��G
o�G3��nFS+4P�"�(Y.���Ė�C|�u��vGW*�rGS�C�ً���F�v5NY�=����t�=��
,f�R��� ���Nxv27`+�y��"��o�P�
���HǤz&�f!]'S��>ajv�$�4/��#�	,�y��[���hVP�7
>�iV�q<]�R'0e��K�$��f���w��_��FV��x��r�(Lj%����!E�/?=,�9PhY�S����;0P��������1s�=�Lv�T2�o^��h�I>p��ٲ���7��-��
Lm�h��S,�9��=��s�Iɖv�� ���jͪ��M�:s���*�B6�'y��W��o�K���p�
���$�`\i�ؗ�����A���t�>���$�v�m���������*�y?�A0��	�do	�J�>�|[���� ����}!�{���&��'�z;�$*��~֋-��hn���&��y�����>8ѻMC@� n����� ��ӁLL冞7�y���@J��3�T�ߔy��O�S��
Y���Ʈ05�J�ɀ�n�:e��qH�����:w�zp��G��w~�҄����|Gf��] {�<�U�7�45	,Fӣ��#N���2���������"g�R�ru��n��E6��m 5Q��%;h�9n,6H��fƩ�j�ۑ��v�Uճ�#�v�+�Hݓ`$�	�Ǚ7P।���vw\�Xr�-�)�=59���Ȼ9�Id�	����Z�˺�����^ as �nMIkkSrVx�x��(�y}QFo�j<ﶽA&���Ju�$S�����7����۰��A��2�/��pw_S�@=Mk^���5���2eT�}��@����:,��,�zc}��	�f�f�T/ܿ^a���r4I��|s��T��?]8~��el��S���p\hp���;�r��߰*�r6F��,e��7-�v�ڤ~�ԃ�����2�WݴZ���\_�l�/�p��-m�a��)�5�7��ؼ����F��w��j�d�U=�*��Ab���;��Z�	b�ύxÜ�~<B"�sRs_
�T�����}пhjj��3�?W^ic1��wu�^��&��S�����O���ah��ە�:��U;h�x����nFnU�e������߾�$�|��4	#���!��M.�����i���Z%�
��>O\�D޸#K�&3��t�%P���k�=M�Q�����Zѱ_܄�Bg�CC}��|��|�T ���,�F�������X��)Yn��f���`j��a���v�_غ�� lJ�� �WG_�,���� ���Y��3�TDn�t	6|ߙ�l�mْeҶ��x��G���WU/���<Q���������2@F�(��y���r�ߢ�Ҏ˳�o(4�g��!����¢%]�Ȱ�1^��1��⧟�p��)m@]�����ѵNlQ�����\=X� �8ؒ ���<R=T;��"�ˬĘHXM����5R�3��¡��@Y�i�NM޳�SZ����D��j��S��I���(��1<��C��[��v�+��"tL���
�u���F�(�m̻_z�Qc�a�^m�L.ΰԶN�~u/��,^bĂ*�4Ψ��oI�RG,�����{���Hr�dhr��u'$��p)+4�P�%��jz��9�&�S�!���XA�Ʃ��D�|��}E(#�{*e�}B�^�e)wE��ƺ9DS����)-:�/��6Q(+&��i�'"ۍ	/��
�F6
Q ̟M�a���C'T�F,�q�Igp����~�S�[��M�@x��{~�Ł�mrs��J@�g#h�CW8�O{��j��&��r��*�����ޢCó�/߀Y�{ȼd�J�qc�Oc���w�4��u*J�����n�a��!�A~�z�Qt}"Yf��;Q�PD���j��c�	��p�:z�vW��)��J�|a�=r����,���tm�E��?X�ykO��*u0ʡ�F^�<2�}bAw`�#�E�Y;5����сQ���R��g�9�}{�U4`��$��������Kv�|�:�s�$s�Χ�ۤ��Y�֣��:�ڰ+�_��gX�Q� ��T�J���I}D��᯶�9���H\�ѵƄ[�N�^+@�V3�&���ƙ���*ճܫT�f8� V�i���Ov�Z�z�t9�B�`����.LW�>'�
Ŧ|N�M��W�Ķ��>�4~ɝ�=@>��Fi'*$���c���:�w�p�%�7&j��8�(Oh���/�:18�!z�:��a<��0>�;�a�#!�WU��P�?2������r�i]���n��`��K���"������>�<5q���#x��L��f�y��A(�=���"�������P0�	��\\\�}�ƚ�p7��$�)2�r�[Ը���~a;M���B�� 9����S-��Wu�ce�s;�O��o0���kM���/l��Z��G�_Ù�K0����X̥�i��[H0��Cg�H�AN�q۷U�n\)0@ ΄�7řs��k��өw�6�9�c ���lpն�`�_�W�b�G��	��;����
�*ݑ�����Y��?'�a��Q��-��J����	?vLC+�-�_mb;a����JD|������S�a����c����ή��M{���������oiM~�H�%���"Q�Q�Y�(s��.�G�G>�)��ڶ9"�4;�>FCX�i]���2[��A�5�@�~����v�2z�2��Zc \�	+)�E�����C��of��A�b��f��)c%@��S�1+הoy̶�RrYe�������V��5����{PO&���Ʃ�E�C x�W�G-T핧��f��c�� 6z�qb��9IG��yR[�Gx&�@���<ׯ쬬�.��/)�����3�2C���������, �����	)�������\�Ww��>��Ԋ$�u��Fc���P��������u�V.�e7.��.�-����u-c�42��H��k���X�:�;� @g$R\����L�����ӭ��C����W�a��N�j^�^!Qv�V8�G���L��e�����m�x9��9��Ф�0뇆�d�P�ƈ�F��8��!V)__apѯ��)����mo�W"߸#4�(�>���]�f�����ݚZ����Y>E�
/��xӇo�� ��y���2��\�^����_�8��	���C���qK�%j�*0��P�U^f�`��n��5z��4�_}�snఞd�����乆ŢW�)�q�c���AN���33`C�X��/=.]t���.����y�����f?��LB��x�c#ݧ�z�#��������R?;�N4���Y��'��EO���%�+\wt~8���JD��~ʢRw�4F#9U��C�Vֿ=�����s����5،߆Vz0P���R1T�n1!v�6Xʈ����}فkL[�bCE �ρZ��Fvph��`����1���9(`UJ��"��W
8b�:o}���%����W6��?�H�`f�b)	&t�ϟ����P�j�&,�Y	|���+q��S*zp�kʟ��6G�Z	fA��y���+�4F	f��ψϚ+�j��|���Ls��IV,Sk��e�͎S�ڠ��s+ͣ�v��ب������Z���2�h�-- 惫dV���#�fdv�b��X��y��i�VW�J�ѯ^��c�N�p�c�2���ee4�լz(^�va�D��ED�i��Ӵt�/B�:]{V���y�eo��z8T�-�L��=G��B�@>��s3�>�љ���-�[�7�(^zv��G�x��h��,:�pg�Ý��/7�Fo�;l<�@��B��E��tw� ��Q`�7�~��l�4�4 8y:�i����2C[��V.Wٚˋǣ���o�!�� C���=6�u��#��ы������֒�)�J�]��ޘf\��"F�Q.�v�.w�2w�:�9�:[yMg5O��k�- ������L�.��B'�Ee�h �2ddc�	F�g��������z1�Ü�]��5N:����`c$��"	Wp2�k�}&�I�.&칺���6U���T�w�"�w�`y�AI:�t�[y��� H��ҽ��m�=���e�Ne�v̿����j��)�,�B6�(��&i�5���$�k̦g}�)�>�Z�%��������.��!�'�Z۹�$#?��s��do��'0p�%���;��c">EfJHs��̏�>LYJ�~�d�h�ńjIA�s���� ʬ��\�*l��3�_�K�mc�<ۤ��D��o?g�cr)m�[�!XM��\2�	d�DH�jR?'�
'i4�=`q�Ͷ�
�s�}�4��`D|��x�����}���'z�H�(���C /HĽz�q��g�¬w�~ܧh�N�k ���]��
O1�`�Ʀ����IզQ�L�c�=��X��'�{��v8�O@8��S�5�\j��Lį����!_�������'+�C[�Ow��a�'yu���Rqu���u�4D�Y� � �c
� ������1c�L��6��u���sjk	떼�K�/߃�j�Zn����|eq^�;i08bƀm��#TUT�\�����*�O�\�'I�	ͺ����c��1��r!0,���!�N���� � mD�����|�����M�g������E�������`S��v�Ě�x����E�8X�)8��łEٹU.����� c(w�RۇXYY�M�譕* �JIS����XB��k4�T'd8h��`���o~�?̸��CJ��W�_Z(E�E	���Xc���e޺yI���r�B*�?G�J���^�t�*יY�R��Z�F�V=���r�d/j-p�]��{\S���1�1�+�xNo�Mw*�"#��.H��C\\��>4T%MR��YF���R�s�Yp�:��VU�Ȓp[dVT�i�t0�56C��m�
������������y�ݻ�Vm��FmI�.ڷr~<3��d��ъ�X���B^|w/����#~��]6�U���>��qܗ��KZx2��@����c�jw���޵���{�YX̝��%b��x�i�p1?�-��^��3�Q_*��)������CJ��\.���`�w�@
������Z/�An"z���qhA�|�7Yk<�Y���q�k�|�S�ԔyUl�J��l ��M�ܲ~�ᯡ�~ĕ�����_ ��
��p @������x�Wǉ`�L ��y����(cɣ�&�+kmބݰE�8D�@ԀLƾ�o<H���pꇅ�b����$�M4����|�ڛ��3F_�I�YY�{�%�66��Η���s���opr�~�]���1�<���#�� ;"Xx������H�R�:�����F$��c�/���..z_�D���`펃(7\���VWCEL*3B88$��!~�_&� ��_�c�� ���!܄�KRYY]�g?X�����)u�p�/sZ���a�������9_E$��PL$di�K�`��é�R��U�\Cq� ���^��śƯ�5��{�F$|u�5Ҍ�NL����ӝ�:愎�%�I�DYݔ_��p�<�lŌY�������\�u;�`
ͥ��(۷��&�|�)��]f�{c9�{oBB�Z���f�:��_�٤~}�����d�F��;[a�t��
���P���r� ��	�-�9�?����=c�W:��(L͗n���մ�3�\���tG���ś`3�E,~VL �'�;gg���d<żԵv�JT4���+��u����R�>���!��#_���;;��&0���5a�����\p$���̀����<`�9�^�D��s��z�:A=��,�e�������%64�V�)S��|/�Q��x�b��`���9��5�Yi'\m�-:���U������1��］n�	l�	Zb��&�du��������dfE5��+x�Ӆ[�H�g��������(��La�u�:��=�噧����4ع�׻�����C(
6�O#Y�����bu����HD1���>=�Y���`-�������!~S����:�S�%�@��&��2E"6��Y1���5�5�ru����v$z�u7�[�rMCAa�-��2��R[Gmt튞+�z��4q��	�E$q�HM�L�O���Z���#�����T�T�~��]��;����`"x$��z��1�nُp@��ݘ��%��444���9����F��� �ɮ!����n��8���0�Uɰ�]��������h��}������U!����K6��~k�9����S�2B��e��P��£�����:U<��N������Jy�����|��-"��F*�|��"YΊ�t!���t�������*M>X�\�i�g��"�����/ɴFs����0�9��n�'+a���L	��v�t������j���񜷝���s����{6v6��oz��L0wW�^u[����S>��c��h��Y�s�����~P��Yu����9%���6�Y�l�<�g�膳.F)��i-j�Z1��eyL� ���@M*Y� �~:S丠�Q%����]
�J�R�Cӧ�0�N�l����ޡW�����E�CBB��'��g#BG�Tu_���W)��ފ���%i��
/V�^�ޅiW8οw�&'}h�"ߖ��Н�2��?n��GC�y��Jl��*�`W���v��#��ga� �C=��ټ�/H]��P����|�����^���B�W�g/�D�G}Ԩ�H^͊��L`Xg˹@��T����z)� r00��a��J|��%i�2�lx�j��E`�^{l1��}����ډ1�ܜ����YS>]�������d�z�Cp̥ d�RD;	6�a`eE��>��xF4��]=�$Ur �z���v���#��H �Y	j����^�?%��)����;����?L�K�Z�5��Ϯ��d��	����G��� i���$����WR�	:�3cp%b!}K簅��!2�g�Æ�/y�_�P��8R!?'O���F�k�����}�h�&n�������*Ҡ"���`��PJ�|y�E������ŝ="BB�'�]|%�# ���3����o���-��D�\���a��/�)�[)�كM0>hu�O_*V�ǻ�Jt�����_m!�f�Q�u���:J��NR�����\�1K��	Y���Zz�A��:��9޿`�Ͷ;� V�U5�Q�U���¤!��ώL&)�]�6��=}�X'��=m��qpWtr��4Nk=+�0�N�C+�iŬ3��AX�3��ҹ��og*DQ�h�;�=�������C C�A-�`4��*>'ܿ�p#�;�$	�M����+b��lJP#�N�������sC[�\�xv5�([K^f��%����9�Yx�F��븂_���܇Wh^T,������ld��`�3^�,%,��sٰa�����UI��pX������S���t,����H��B�H˽/���P���) ��N!���LW��0���O����i��Ɯ�>L,w�-�ʈ�p?�<EQr$nG���{ɘ�;��^mŮQ
(�X/�����+' ���M��Q�������لs�>��憎���tn��:k]�4��/���>�YEƮWI�^C�\�R��Jv$[�4�A��ݥ	�=�J��R��S���ڷ�t9$^9����c����B��G[CF3� v�T��l(.ao}4��P�G)�����J�8�u�]�����F��,�aL�<��>�{@yy-0�:%�@�P<�B������agAb�V��$*����C&�9q�YrY2W�Ϛ?^y�s����x�(@�ܑ�]���?r2��B̥3�`WOs�goD5���bs��<&�>��R�pP�2Pe�G����pG�純���.=�_kZ�^�D�@/S�Ⱦ���g�{��o��s��B���ÒBh�������֒Ȗ���@̂_:}�: -�$�A)�o�VE/E'`��Di(T��2��ϯw`KhUmm*O�������ꛜU�D�g�ӈ�t3�(<�P��r���+�D �y��b�Z �7�z2�K�+l4�@���i�+���%�+Z'��EG�f���P��o�h =��&��Y�'�ޓ��$�q��fv���2��,�	�39�ً˨�
���ٚ=�,:{a���������:�����
x9 =u�+����D�"�X"e������[ߩ���t�����n�+�p:x�wA�dy��ј��e[S�M"���8>s�Iz�&���ύq�ɳ�2�3�!�g����[+	�yN�+���xů�#�������ƻ[�(�{�^�.$��/^�_�xE��pN�f�U����+��{�z�)�M���u���S��V<�*|I
;������H���'hmO�=�r�����$�޷�ς��qO�t��J{Ӎg?x�����9����s1��0�LT}��R���~7ˍ�~��������	N��8x�2=N����<�<�p>k�)�S(-!q9#�<�׺��m�hB�c���g��*Kt�,�?��ͳ�E�Me�뤧H�M�3,�hͭ�=ؘ�,(�}�[ׄ�ܪdD���oKן��r
D��5��
5=H��Q�ӋN�[�d��N��@�����d�y�ls1v�����|��b��ڢ>�
s7�q�|�;�3Ɠ��'��i-5�$>��j����=���$t�_���l���Nͥ���b��}�1f��4/�*	��ċ��\=7_*�GXf8�bd�~9��Do����^��a�yL�����d�'�MH6�j��H;8g U&���BZ������L�O�D�zZE��{������q�G��$R�2u���Z\��Ŧ* �"!$)9ހ--8�|�z��({��b9����Ho���̍G�箳�
��)��~��fs��_[��@�t%ɷv�рQ)����	��h$WJ<+=K�C_�x�0[�j�%��<\�<�z�?�-Rͺ��]R��
�?���]��*�2�繽���m��*�)2z����+8���`=N���3�!�*�A�1l��\��8)|2ff�pвяK%u[���E�R��g���%nˡN�e6��勌��X���ݕ�8%JP�!s�|k��}���78��Y�=f�4>CI�	J��&�7э�J��P��<������4�D�Nn^5�Ҁ$�fK����"A�{�lM�/H��Ӟ�.����;;�`�*�QSX�8|��W���1�%0Yzrj�`�����"�B"�fS蟃�5�J��!r���53"}�4FV.M˅�%�`�fJ	�L1zP'�V�Sa��wVdUy.���7�0�'�Qؔo�\�bM�i'_��we���8��;two�T{�����5:�z\^=�#��=�Qs�S떔��
]#�>U~"��o��P?�]��Ib=�������m�X6���pa~�c[`#��h�&�t4_����ؐ�#)>�C/>�,r�?��/�	24Kw��� �0�d��Ƞ�
��.�&�^ҕ�PY�(�����Md�%��%y�eލ3FM#9{������ub�ux�%�!����ӹ�0��_�T������A������ظQ�Ŝfm��jv?^���f�,�^X��I,~ej��:��f]0�l�����>��-�}螝�ǒ��V�f����`e����E�Z��ʢ�k�#���b��F?q����@x��j���Wc��,]�ćüۼ�>�d���`IWt5�Ftn�y2%���[0�_�}g��h�-r��V�F�8�e){2H����*��.j�9z؂~�K�̞�����rd]�oo�"��qNξ=ݑ��I�v��~c��p���?��I)��πW��������:1�����A��5�A����������yoC��UTk�".��x�X�uf>�;#[F�k�g�v �ԕ7�?���ɰ$��t�EJ�����R�R�0B�� D	�1�Fb��ݽь�{������������u]��,r�c�-to�r`�-�+��%K��������׆nC��[ ��3JKKw�^0�e�>8	����tIC��U.iI�)0w�W�y%as����L�#O�,�,��H)6��R�sϫR*�G��;Wcuԅ��u/,�E�ȴ����Y&�;}���I��_w
w��g}u{/t�c�I�Ȁ�(���>&|`x:h�.f��Y�~w����?"l�v�qMj���.�s���R=.��p��U� �Ŝ�r*�(����;�Hoz�9�O��z_FkT�*Ro4�ғ���"�����P%��D{�l�E�A��E��" =i(o��&�ZN<`}Z���Ģ�&�����\�L遆&œ�<GE%W�e����%V�t׷o��t�/	�N�H~z�*�=�c�;��#������MлW�5{��7�����4��d�"g�O��� �3�*�t�h�+����Xzϖ����1���37�U?Z!7���.Z\H�{x�-�d����Qū��/`0���isoo�L��&��aMq�E�`uN‏����Մ��H�5ت�ŹʞF�l�h���[	�NC�(�d��P�%�~��o�$��ݽ�z���6������}��ʸ�n�\Oi�1U�5��/D���Q}X�B��2d2�E�΅��0+��.����j�������ܥ���v���q����X�����Ǜ|$qM- �'q܇�s�ta�u�'2p�Wz#7�Le��RUh���]Y)�(D��v���c[.aI��w���}f��`�7�z3p	����0�g�oD�&�0?��[J*BI
��IL�Tz5y�qC.s�颤�_�R�y��.��%��W�am�Gv��ҵ���~c��X�&G���+�{Q���c���ez8�ˎ�^[��+���1�!ɪ��h����Î� j�G�g��su�n74x���ޭ�!����l��/3fbǇ���J�tc�#-����t{ܟU�#���ٿ$e�\#���mk����rǙgEz��qD��;�OOBW�쭣7X+��dUg9��f&%�SX_�A�`���8 ;�)K���ȁ�<Wuou}O��H�z�.
5�a;o�̳�����BĦ5^S&K��nv$��h\��3�2.�NZ띒�("d��U�_/Y�����8ռ=���8�,�L�kE��&������N����t��kGG��P�W�D<o<��s�Vrk�[1^{���w~���>'�]����C�벨5�o#+��Sb�]�8�MCzl��	��i�V�k�����'+���K������9��3������WP|�&��/�땝gr]���`�[;�$;gfԸ�_���`�lR��=�FG����d�5�|9��֑ˇ� �ѹL�(�����#^k�߀�L��|$se"A0�$��=c\C~�uuą��1��ٙS�Z�/�M����rs"?�K�h���%��I��s�I�S�%��B��<j��N�AIV�E�[z�����Z�������"�;B�	dweq�|w�D��9پ�ЋYX��ż%]�۬x�y)���ꢤƷJL7w��`��{Į��`�� �,�+Y4��YY�gZ�@�T��Zaa!n��~��O����T-����|xX�7���=b�;�ڥ�h�`#�Z*�m��(��`�����N���17p�m!��Q)�q�g� R�㯏,£�ƀ�φ.�!8N0U��	���^(�m��\'�?�P���]c�h�����?\�|B����	g��ͭ�Ƨ��G��b�Ճ�y�Mw�O���y=��0"N�̫��Hk=�~]ҩ������I�;t,�cҫ�M���JiB&��H;�̕����`�a���"y�ƣg#g�k��1}�

�W�7�;ӎ��Y�͕�~0 �;��Yd��&⻯p�R��5�pq0Ѕ#^			��IW���L%��{E��z}B�.<B���cPd"C����������sq�@�9� �?T淰��b����Vt�+>K i��ȧT^���?�*+�/s�ژ��L�e)Yb9�苣�aH���ȣ��|��Pa��s��颣�J�;:v�$���t�DDg0���j;z�L�p͵��p��[���33��
@��Ą^��A�&u�������I�<ݻ����{x�g���I5�B��e��$��Ջ�<�Q���6]iR��`NH��$�J�x�����$����xjtַW��d����|���g��*ǂ4H�5E�Ip�k���ja+��&�k�G��W��`�¿�9��c�ůCD�_@��)�@���m�/ӟ�ݙA�VW�����>fD�����	<��.i퇹-ގ�P�`0X��Lq��K�g�?��R�Q��ǝK����lY�+�R{5v�aL���GHr^>7iP��L)Gb	 .�C�1��="]���:(涓o�>�I~GT���HҶb<�"J����o�:吨�����eP4$*��D��$8��R�<R@^iy�55t8��྅����$	ô7���Y���5�޼y��+nxb"�����p!΃323[��:�+�����M)�<�n�	��v\��R<���^��OK���h���j�:��Vt&��nI�b9���s�ŝ�נ�$�N�i�ެ�<��^����.�}�j:I˾^'N����z/�q0vM��y�(ztgG���$�3��n.;��2�~�vI3��	���C���ԗ%	�W����.�}o���#'�fz9�0Ш��-�ƥ��h[��;k�L���q(z2��8Z�����(u�!@ѵ�`�čj�ێ�6.?�50��b��,��uu�JD���<&��}�=��ZP���mm/z�i�����O�3N�H�`�L�݁�����	 4А���>�䥆�a�m9-P�M�+�oo�#���ԯ�)�m9b$Z��hgq���]�&)��܍g��y�O*���%s"�6�2u�a[ �a�.ۏ�e�Ɉ�������7!��s�Dh��N{��?1�[�YK��ޙ��$]dX'\�U��>�t����ר}���&tf�S�<�{�|Ձi4�L�����j9Qa�x���bp���YJ#��[�28;u��ݩ�� j����ׇ]��eŅoޜ�p͆m]c�N�'ai1I[ާRcK��� �^�����0V�L�{IZ>�q:jq]W�q�}�����N]��>�q�]
��fQ��M)ymM����.�CW��xYK�{k��^,��Y��K�}��`�����QʂH�D�����x�e	�����Prֻ�qI" S.)��>9.�Uۍe�����2�\��>p�P~\z?P4 ���t���� ��u#3�9��7�prb�G��AZ�_������H�?�?�4f��Ru�"��f��Y���￞���%$K/'���3�N3�/P�]�{�s���涤')�q��x	^��c����'}Ώ i�m�N.�,��@��A�Z�Ό35�m�[�]H�$G�r�X�0���TyE�����#1^��z$�~�ߣZT�٘�O�����G��ЯJ	0�@;�K��dK����#�&�Y�M�F��.j7n�_��P�PI�
O}{m��h<	�>�n<u����
zg�@C0}���Ks�(z����ZѪ�.&�߷�4�����3]��hd�h�k?��@�{_���ge���(�Q~��`�ԗ:s�e�C���@�
�6�_��J�i��񙮁4�������M�<�B��Q���#�p@�Їyܔ
 �Ē3Jb����H�ƞ%�5<<<��"���Pk��8J�^mRz��0"e?�J$ć��$�MEM��LD^��V�lv)�f3��V��fj�K�#p�����i}�jG��.��t�=
D�
���K���������)sF&��ϳh��^���~q�	���3����q�}�p�@[�UPPPf����\������D���o200�ʔ-3�"'�������P���p>�%M///�7TUU}��0j���e��N'|ϡ��d��¿�[�1}���@��v	����o2�=ԕ$g�ţ����gᄑ�R;���o^{�$�v%��T�DJ���6�}h8����:��7�<��؈�8�v Pꅖ�FP��钮*E>�:ύ��k��8���~��pV�Wӵ��ܱ��S�Ò��ܚ����S_�p�|[��2��/�Y����G��{���y2kx��xb����)���iӢ�������L��4�͑ۖ�7�~h�l�"�///ŝ�_d��>q�	��]����jҙ��j[Z�#X��-w�T�ۀ�&��s��"{�Do���m�Je����JU������օ|%��/r����WC^;�.�J K(��+���%����Jl��)1��������_q|zKy�Z��'nó�jl2w|w��<�,���-ǋ�b���&� �}�u��}y���c#���<��av������� �.v���ϴ�~�W~q0S>���=����k'c��߿_c�D��`Z<�Ԙ5�#q?��\snn�n`	s��n`svrx|���G�D"u��%lmm���ɳb
׃xĪ�	��u����(%��=�5�H�7U͒��˃�rv:����4Kpp(�$�����	��A�@3յ����O��@`ӕn� ��w;/�d�O�v��B�N���"�@��>~��bꍓ�#K���]K�=�w�b��}~V�ꥡ���^&4�pt�殕�nx�a��OW��:ʯ�:�$��2������i��g�d�,�>�e�b}���;���̶iY�J�^�-�
oy�!���e>�ܫ�v�9߳<��$�`k�V�?8�w��s�,���џ�'l�Q����?[���s�����{yM�	jW��d��R� �'���f�.����_��W���Z�5�\��OZ�����L�,�{�\�$y>0z��+x�ɪ���v��������`��`Y������S�5�ĚKK�(��R��{�G���3�v�:��`��7وSb��e!w�Z�V���O�{�lư[�沣���+d5��t�����/8H4v��T�E�	�+����/<rv騛D��mq����$8������ۑ􂝋�C33�11�m{��S���Z-�%j���⚛5�_�{xT���<�Y4ܫC�(P� YH6c��{�~k�.�����`#"���w�x�zw&�**�lS�o &�Iy�[�?���%{]u�r�j7j����q���-��y�񍏖�������%�&o16��Ck}@^�O;3���>��/@q�$	iA;�k����������4�ާ q��n3T¦��ۋ��$S��b�K����̪W�TGB�2�v,��oz��-�S�.=�?������H0j������O��Ĭ��s�]�㝹�o�W�n�R�؄� ǈ�zp� ���Q.����3��E����rvB��/-�����M��)©Ԇ����}r�>�'8��t%GI@�2ܒ�V��CR���ٷ��A�+�6�"�(1@|����|�����O��� q�ж���iFpI���0(�9=�?�  ���!�j�`�,R^4��``b��?Qe�^ڙ�}������]�
��(���744�y��TUW;��R%x�O������d���PܒK�^RcP?��6��h�Dk���Vdb~�q��է6��6a�h��K(dٲP�x��A?����r�OS���(]_޸8�����K��DoT����l�E*���gu>�7Rڝ!�b��X����~�䄿tO>X3=����f)��v��ɹA��˙��=�t�b�c���[�c��D��D}m��V ;�r����iX�e�g؍���##�DXn,9������D���c7ww�Ǝ��[�����C��(z����/Y{�8�=m7��f�%��wܧ�@OϚvy_,貾���릲�J�RZ�{��W�KE/�뿲����G�P<etv��$��fb�V1}(���m�R �:�L	kF9[ x5�b��psE��0��.�ʍ1�ض1Qx��!�w���܋�����q/�-1�c���9{�"��������2�&qO)f�=��S�\�<�"��m��	B�pw��XYYu�l�V���t��j$��)��cr��~Lf�s��-ҕ7����K3�Þi�!h��RE�Q��H��l7:��-���Zk
_�/�����>�Ը���A������y#���Y=�}���1��B$��鄹�L��lI �'#`�ORMԍ�
J�a�ʂ���vn��vJ�F���$��J�K��/3n��֦!��J�ɣA��$�~g��㿍@y��<��Q�7�p�5!RL��7��X�Tp�׫�|�Q�n`��ϧ�[����Ɲ��P�����v�8��W9�T(3-����m\0�OT$����r�����K.'��$?����%8�����/��Tˤ��R8�-�4�9&���o�6��A{�U�S}���T��W�0�2��N����r�O�s�_���P����^!G�?�݈�t��iQ��,�Ey�
jx0�2\i�"F!���l���/]��`��#&-��`ebaA����'��q�yW���qW,�Z�Y GFn�-��Fσ��!�`���ũ����vv|	�z55O_}n7�Y�5ITΘٹ��,�y���@�l;ۧ7�o�h��l�Ȓh9�啙k��څ�q����7�7m:#Ѻ���3��Aj�H�����uC�b!'Atx}xQ���؎�]΅��eex�MG���`�38]�iv#"u�~㾔�4_�m�X���w��[���3'V�u�O��D�3�eƿ�9$sM4kx2 4F�\�>"�pF9�x�������<j��[Y��<�Fb'��Y�4�P�#����{�cc: ��a�Y�ō@2�����w	���Qs��xx��)4��aܠP���`܍'��^-f)F�9-�YI��2 ���!�s����A��98&^�j�v�3��T,�\�vy�f�[��o@��_�y�$�(��з�]k�rB���G�g�dսl�z�an��;���x�4� Z��Ms��x*�V|�썄W�/�ˌ[�5���<�{��%j�fP�?MG�v���N�bbGǗ���^p������PiR�--�)�>LKKK��c���N����)�� j�����wB}q~I�K8\R��`���9d}=#n��ή���`hr�g;9cn`� ���pD�� ��)�J�,u������S�V�Y�VR(~gu'���W%���@K��$�y����M*�?W"�g�+�*�\"6^�Y��{.m���ʟ���fLN��b<*���o��d~M�3�p�9�����o�]��L��]p=|��K�ϴ*N�~϶�<Y���7~�$�:�~V�R?;?�j`Pbrx}!�E�&��oT��s�1���0������UT/��N�x������ַ����Xs''ʶ�6V֎�Aʐ��<EvI(555�G
4�������H���4�'aU
�RK �����ݖ���=�}�N4ų~��Na6�q#v1�v�[�zҜ�u�����S�')XR����z���r��3ukx8Ť�o(��Փ8Y#zH�ɝ��wz p.���[�1��B~+A���A�Y��3����zw㿽5H�,���������cL��fmW+�{VP�8Vvv�BQ=N5O���\��֖��߿I�ɭ��4�]]��{{�m����o��wW�_;N�7���������L��C��agg^O�<� �ITT��h[;;܏FGG�lRG�g6}e��I[t�=���S��u��|�� �A<|�4&`�nM~^>�Nà)�v�/j��04u��\:!�t����Wo�6���9����!xyZW@7���֍���b��RC�&ҹ�V4���3av�� ��s/��1~���Pwd"RT�_�u�Ay�q_���,Z�����rb�9�R����w~���n���X�	uf'��f��.��/��U�����l��{�����}a`g�g���5��͍&;;����p	?y��9a�|�㮤��p>|4!�XvNNμTMUUFv���������I�0k����W�2{Bb���5�C�w��\�C����Ip#�dP�)��������27��I���Q����i8a���%�,�Ʃ�dt���B��`|{o����ob9��>����Ǔj�I*��A�M�J��� ��Y��Z�}�j�2�_�6A�w�5/A�Z��.�`����������{��k� |��1�������T����x.�e���=3�}�n�ck������^����6�mn���S� ��/3\�q�>L[v�ل61���5��ÏO���y��B����&I4����o�����Mݐs�M�`�_�:�B��~����eT�;^�%W�}-x���0������L~�N���rCc���L���b�.Z���^��b��M?j�L}�M� }l�p����F	�c���)�|��H�Ph�8Qm���	��{��g�R���L7�O���̓;u�� ����[  �����(���v��	���\�4I����V��%t[�z�Rzy�൜��ȝp ���L}|� �V��)�231��T����K�|O��n����2X�gb�R�hV��*�1ڦЃ���TZ[k��ϖ�f���b].�Y��$���I�D���'�4%r��:OF�����GY�UR�����(7��#Z���xCf�[i2�D�^!Dhy]祊2�q�@R�0���ev��v�M��x�� "4ѧ_�wc߽�"XV��Q>�9؉Vg�Y��K�r��օȿ=�+䙠n��3���h�g z<"����-Ƈ��ڰ)�*�1b��{�6bNuk2h�ޥĜ��1�I.�.@�2[�/�17�eB���S"Ω�Z�n�;�H�آ+����W��X�U��eF����+.Z�*ff��6̍T�ۅ�$�)��cܑS{��r�i�;)��y�3�Ky����BwG�����#�i�2�Cp�i� ^�\oU�r�q(�K3E{�n�?�����"�G#s��.
�g��;�
�� S�h�mV��5�ev/v�)�eP����hR���ڃ��Q��-��gRN���G��M8��Y/qGrWGYڋ����Q���iVaֱ4����^C2ˎ��A�*��"�Ww�2��-up����,L�u0+!!x�z��B��-z�^o�*4�r�R'�9o����D�g�怯�*�}�i&��[�ۄ�\�o��������3�z	ѭ_U�M�Tl���Op��F��^Z�����LU�u�5\��_,H\,St\2�d��t8�Y!�<���3����/�������~<�?���D^�Er�d0�C�h���}��o86-_SJ(W3�0������z2�f�
�R�L��c�� KjJ�w�C�EWz^g��-K�t`k���X�N�����d G����}��"��ڦT ��?]��#�+s]��Ƥ8L��#6
��'��p{)�ݎ�j�v�]��b
3)�V�O6G���O��ud8�<���gb���fa)kM���R;�mq����-�Q8�Ӕc�>d���f��a�(�I�Zv�c�^�<`���큺�W��N�Y�2Vo#��V���뭊�3��
=	?�O����a���:ϢP��y�E�.Õ�8t�>�;��1�{�-k����-6�cAq����򞎕m�*����l��Z�Ɯf�Ŷ��!x݃G�UA(��;n�"AC�����Ût��u�"3%İ�����/�'+��j[^���&��%�]��4�����^Dl�r~Uo�r�-d��)Q�����bgI��I�1�چq�g�i/���E+nK��W_ �@ɢ�̴�z� Y�}��	��n(��=��E�%rn4L�������Փ��f�.�0�G_�8���?��O>}~1Fr9v���~��A<w#=�<�l̲�݂
�9�ŐQ�a	�tzAE�x�6G�u7L	�<��o�4N�z�9k�� �Bf+k� uիUk��z�Ս��瘸��׫eKH̦?��Y>�O��c�/BpGŠIak�w>)������8b��Χ�?��ç��� ���6	a��;4YZ���ְ�ٴ������}n��EpT��R����8(u�
���<���,��Z��`����Tʇ���9��nJ��I�C>��x.�{�*�,��8�W��X$��ίmV�#Pv��c�C��z\M�5�@f�{��\ʓdr.r?�%�U��#O�����-�6�OzRT]�&�-�i�+��O�(w���vA��z�K����[����碌��I�'�Y��Fr�-�W��[1ϳ�SM�GjȦ<��̈́s�A�"�l
4K�1���S�֒�fFj[�+l���I��R��Ty6���{e��|��3�e3��-��T%�������7<3��Ŗ&o�������>'2;���
ӱ��n#Kg*���3*�kv6��E�RyWy)G]�Rj6K�Fސxh?0���?{�JҰ%�`r|�2~�lNX��G�Z��$R�i���g��ih�0d�ȓ���IOy���0M�q�F�����eȆ\&� {ɗ�ٷ�j#��p6���0w�Mn�#�z�&!�:����,
�G�;�T��_� X��i�톇QϚ�.�@p� �8|���,�Z�v=���C�St]��. ݀]�|7F(�ܣ<�2�/ ���2���w���6�Q�܉{��Ơ��g�=ρe�<d�f�,�Na�.�\J\��4�s�|I&p2��]_EQC���1E�*�����]��EIt���I�QB���i�M�O#��eRj���}
s��>���Z;DJ���0K�(K�E�L��O���\��7�`��\��
I���8�E�=0��	G�w��|kQ����i�y���ʗ
h(��h��İ[�N�@�t	�/XH��.�����h��g�z�`��U��u�$��T�q��3BK��#g�I�`��ƩǂV�)�!q@��ئ���kN��=N�x}�sr)r��K+!���&[/�p�?��6�D�)с�,�M�f�͍U%�( �`�E���+:����`4���B���������%�zUʷW�i��in��D#)N��x�h#�uFk����x8��*ulIg���/�?���� _$�L���w�d�8����S��f&F>'�|>��ǃ;$���?��N&�
drS��~,�i�٩4j�i��o(�������	��*���/�FR����k��0��-Q\Z9+�2��q����!��3];ǵ���pD��U
�7��3�T���E�����X��|��V�W����3����{�H��-�+��tڑ�EfhB���1�D�eW�ƭ'e=gH�qI�?4���>}�}>�n�Uƛ�[�����e����]��/�M�~�����fu��׾h���Y�a���jՇ O��<f�<( X�`�zs��8N!D�,�]��>c���c�����#�b�I!�(��~�C��Q��������$<dUgV�|Wʓ�qH�%��u��GX���}�ϲP�Y�>Gꃝ8����g�4�z_L뼲H���^�x�7`V�o�*Q�!�ؘB/���8 -�nXq�Eg���c�ok/�nSu2ɸ���QC��Ee����&t�&���T%;���>8$�@gAV�=o�Gj��L��g4R*(���=���Q��k��s���u����+�<WǷ캢�袿u��:/��w�A�Ѿw&���s��nCL��޷��L�m���*��P�l�^�����(�)���%����ͬ��e9LT�4ʇpH�}x�'O�u}�e�I��S��Sy�HO��d ߬,���븡j)�}�-&�V7.(�'\�x�N�>٢{8t������k��u�>��X����La�y�RZ��TQ:�A����լ��b�l�r������Ѥҵ��I-���@���K� tAAE������'��M�@ �T��ؚt�R{�9Lk���U8�j��E6G�ף�S�Ҙsa|��C���D���P{��򩓬A�-g�-'���=u�a���}�%y�XϢC��,��s)	d&ݝ\fwYD��c�a2=��Œ#x��%�c<����g����no��ӮE����;ʻ�78���W �Y��a��}�yZ���.Y�^��7A�B�HٱST+�A�QT�1v��{��
��f_�t�Y�M�P�������.S��	yF��D�LH���޷C=��\��:��0M@�f�]ǌ�XD�p��O�@B�I7�r��<u$u��[ʾ���=�>�K���)'w<�#���6�^�cΟ��������Z��?	���F��
�&l�J�ަ��<o��i�aW�Y$�a�Iԍ�%���W[wI�;��j�D��e��V�o�o��C�7+��/��R=�~P)�����^�Za�{����KE�QY�~���l%R�P�H]X�W|�88 �4K�}{}JF�Pʭ�����p}��-6�pm�[s|�e��*j�4"��� �Ir��Ii���	9�)׈�y�M`B.��gq�z&�{����f�;uP�8�=-��"W%�}I��ӛ��s��p!�hST��5�M��Y�w�3�f9D�%�z���{<������'}Hf��|Bغ��=>��R�MN��ǡ�y2�#���+�A� k�	߄`T�)��ל�?���Gi��2\b�^��{l.�S�W{�y���ԑ�Ng��Tz+�,������ץ�Iн3/Rxޠ�q�A����=�����[֕%
|\��ꤝ&N�	7�ڦ�X2�u�o+��U�/�re5����n�i-���v=<�-��j@�Z��$�&�W�4B)�����MtȹG;�e�1���3Zyo��#��$�>�^���<v~pj�&�����_�f
�**�����6�ŭ�W��lF��^<�[z�~�xU��\�c�8=��hz������͒~�p�����&�����7�]�i��zA�l��7S�`g�U��k��,���J�Z��w�	�E[I�|M��[���S
�2WiWg�d5�Z��P���۪���[Sz*�U��l�Sޣ5�$����9P����+��,�2�}�;|���wb�AdIш��S,�m��w��N��-���\���ue<���+w�I�Q{Q�%+]W���A��Qe�w�}�@�8zv=�qjG}���w��V;j���(屖uQ)������������~�"s�ș1�6���"2�Q�{�z�$�[x�I���Gg�3�����+(�l�9i���'�s���xNɎ%�3 }��{�Ǘ�RҬ��5]W�����Yz��Ӽ�q9�=����^"JwE�-�(k�%M��#in��O��!q����q�G_��E7�CXJ��6�f��ϳ�F������vG�L�wţ��Wo�xwPՈu����G�6��p������;y�*��O׽
E!�y fl��و8cN��������N�F�����>}i�WR�JZ��@4��`��xp�C==�`u��g��E�U�Q��N�|�ƅ3ޫ�xl�+`c����x8S/�UEc��9.����� ��H�fg��L�z�!��bh.kBݡQ�/⎣{����;�L<Dm.\�X�XP�#KIZz&| ���9:c����A���&G훫�2^,+X��]f���E���ހξ�N��<Ҷ���^�
�����V_��%�<��^R� 5$�,�O&D>�m�st���Y�%�`t��W�S�P{�cC�|^�Ig���k���?8
���~z�`)���J��W��R ��^l�<����)�5c����M�;fN���/�ܧ"Dw[-�?r@/*|�It@�~G��T_��v�J�4�瞗3c|�1J4�NS�[N��W��hz���_jӱ�u?�rIe���^�6�k��o�9=��j�r�ķSK64ǉS�(P�cu�Q$Z�%ŽTmR鴢2f��K9��?�!��!A���|3Su�dō�w�7�~��oz+��~y�{H�t�<+��C�����-���q$k5�O������][ge���R�Bk|#����
�:IN�쭣��ma�{��!�~VN�Th�~%-0�ƹƴ^7/c��<o�`S+��L@��W�O�P����f1r@4jI��M��E�˸\���7F\��g�s�0%��!n�piK:!�@<�*W�:�2ڲV��Z�Dh�h�G��EhV�m险�?����%������7���CG�|
�j�A,�>���yp����S�p�����.���ڌ��Bi>��C,[����F\z�n$����
W�yD�bIhz�uӵ�ۼ��w{BA	��>׻��� s��5��c����O{��L��b�ڹ w�HRs뇹{�>��1�]'A̛��O��>��=2G]o��]naO��J�ٯ�[��&��pyd���) �.~���.����s��w�˺��e"u�7JRd���������t(;���%��zc��Vn�qd;���p}���$���#M���|)9D���|�u>ҋ���$�ն�)���<i�x�_��-/�R��Y������j�_��>�g�%�u츊a��V�uUg5�hSXDZ�"��̤�����xM@;®�d��\t=���VZ6���b��9��N��/��U/GІ���#W@~��U��z+�2Z���3c��w����`�X�@q?)Y�9%*{�hY��v��+q��>��o�3�ܢR����FW��b�!#�.���꥛�*�>G+�n�~���zf����S"�Ց��ZӛnMu�2�K{���d������0��eS�JOQ��U��e����JG�|B��d�����8�ki#�V��P��/�b�y'�HX
�vq�����������?4�W87�Aj{��'��d�w��ô�;!E'���i�)nЧ�x����m��I��%��s�NR�JV5��!�����ԙ�U3�ɹ[����[�XK��I�h}�@����%��}�6�sz�_�Lc����O;�-�(�.X;�8����9x�z9�ؚ,�2�ݿ�(��ޓ�B������4����P!oE�9�\ٰ��ii�d�������!x����Y�h5C	$b���Ч���8�&��b�p�4/�h/\҃VumNR��IU�K�\.m%�V�����1'��D��I#췜qW�ʵ�j5��/�w��'0k5��E��8zd�Oa��x� ۍg?�yI�"y�u�,���O~VV����`R�,��l��f�f�mo@���"�����l�p���_�|D�[R�4�ɨ��� |Ơ[% ��C�>GP�@=ݖ4�}�n�U_Hq���,��/�e.t�������:D�����d�$�Ąe�q�������[\����}�����k���2Jo�Df�J�ٯ���u\�=�<�����:��:n]�.88ː�8%��M�1�p��(��ϊ�Ua����=ü>����l�J4�i�7�&}�>h2}/����� ����fbd�e���ܡ��r�MHV�[>����[X'D��%��^�e���{��.U�>e��?Dy�p"�2
�B��� d�Fz,���.�TY�<ϸ;�DC���GW_J�čc�>H�Y$�$с�r
{���*P�QA�p���3���L���)����#���g�S,�y�4L�H��&7lO��HV�ũ*q����� �*&6"��$C_��R#�=nHY�}%����uB8�v� �@u������?�tB����ѺAs��f�+��^�HWj�3֏}�r�Q�E+�Dt�p8.s��q�@�c����8���x4�4qwZZ�K������)O�u~��)uL���F������� �]ze�K6���?����lw���e`�V����Њі��t�F�iq�"�_h+����:&��/��j�`ῐ����?I�P)�Պ0^�Rv�� n3X�r��o�ny�!&z��|����M�*�|��m��V�[�q#��|� 1��#���Xc���ms!��h�<>�* �:C^�)S����x7x����/t�KA!��	�(.6���i���ރF�9���ϳ�O���gL7��}�"u�'�[Ѝ�Lb�E�[�k64��?���O�j#����roX��$��o�M�㱯�w��r�H���T%p}bD�VO een������O/Y&�nr��?뎸�D��΅0�{�o�㰬_	U�Ǖ�p�ӄ�R����w�{A�ܶ��)E���jE��j�����x�ӒR�K��6��3p��*��̫�e:��\�[��3��T�bz����[�%����C|íO
�Qϐ�����b0����\2���(Y���<#>�V�8Y$��X��E����N�`�� fy�4u�x�<*��y� �!H�2�ϧ�'�W�����C�N]v)DԮg�ٙ�ѧrSN�QlfI\�"Hy�<�|��G�;����	����ra�-\�����J�S�Zw��;���-��m,xZt�`�3�ɴcJ��]��5lF=(������ʧT�R��������;�ex�
�"GO�Ai֬^�R����R���	�90�и����4���Ad#�P�Km�~ �JfXF��!)(<Uhg��P�L�ڍ�Q�kWŇ���[���N.�v3��\`.Ckn��R�������5C
>߹:0��wT����ϻ�0@�q5���~w���0O�d5��埅��ֺ%���9_���{@8g-O,1nS>sR�>��Ѕ�Ee �P���23}�:�|)��1�нO��h��Y�m}�I�l�`��
��E�Te��~�g�W����ꭣ���7P�iAT�Ni�����n$�A����CAJi�a�B������]��yך�X�����~�}�9�,_|�;vȔ]�ؽ��G�&�t�v��f�V���3^�����v,�r�xo=�-�i��һ��n?���B���B�H����@;�ү.�T�>�O��Ɇ�9�n�K�2f�$W+�*�>�	�fQ\=��R'�(�M�\I��η���v�h�<��Ag0+Zs֔hCXw�1b�?�@n�{�vv� <�y<i��ѺN�"+�!v��r�!���lk�p@��7�Q���E�k�=��ƿ��L@�H3ߌМO��FwH���^R��CN�#nn"�%wt�=����o@�-����}�k[�o5>�<���?|^^��H|��ap+�!K��2m҆�y�d�~M�Ē��+Ih�.d&��<��7���+�c�b���?G��]�
.���:��u�3�s�K3��q�dd$4]I���ϋo^=듹��}Hf�Y���?���H_ϗI"j�����`@Tc��񈅘3�M$�m�1��=���! �a@�u	f{��G�]�
R���}96���i���sQ B(���\�߈�LC��w0�7�u
 i�V��\�+�8mw:���揣�|�Ԟ��bXh!���k�=V�O�9���V��k�v�e����-�I���(Y��>6���,A���F^�����C��!���R�����'���'#�W�"+�ْ���b\�}$��d������VH���~S�b����iFş�4�h��Ӗd٣�69���.�gu��Z��D�ц��,�=�jrw��.��]cL��u4eY.�[�D4���K�+8`��wI����4ŉ�Y^�.�s���$
�K��o��}û�=?	a����50����"�
���$�!�����f��K�l�?�IВMm��F
��?���4�t��Z�-�d��.lP��{�ȖT4dg��{y�3������v�����o����R`�L&�˗R����/u$fj��-����Jɯ[�u�7�i� ����g��͡7Gh��.l��A�������߲�����Y#���S����(�����`d�-[�j�Nڑ�t'.��Vҹ������)qj�����pw1+�3���z�	΅��Byl��~���3\%qEw}��G���(���,Um-r>��BH��P&d�2����@�����8]��J����S���lw�/ڎ��H`�˳�^F���׆����������}�7j.�R�H���a����L	�vr�k��Jf��EJ�̱LŲMN�rjcz���)���. [��d���^R�K5�6ms��W�Mڴ����D��~�jmB7��(kBA��?�K`��a3�o� ��bC�L;���ܒ`�t��E����0�]D�n��}�{4� 7�#�a��ɩ%�T�!��!5�Pk�1"���)h����C�pZ^�Ʌ��p���d�OV'n��5ǋ�xOM^秵&��&���u�����X@�u�sg�>M�A`u������&�X]7�������I��r��U(�y����8-9�Qf�4<��-4�V�=��L)�%�]�xQw�H���i>�I��y�Ö%�$�W�u� ����`���
�����8y�{Q���҃U��<�̘;��sꁟG�tZѿ�����O��;6�0ި� !�;�wH�<�m4��.֬��nˣכ2~Jg`Y��@�ö
Kx���ϕ@�W:-�9U�{�1���_V�:��^КA?�j�=��$�/�1n��K��3oAZ*�QX�\�������/���J�����}��t
p*O�&�ҩ'���!0���H�ےc+8�NI�����;V�ms(F�S�r�R
h�m�zR�!H���~��ZJO���>�� �ݺ��Gǵ"��lgK�H~(������(���x�Gw��A����!�1J�sD��3j��IҬ߬�Q���U���r8O��z�^�{XR���Z���Zh��0��{�#�e����P�6o'	}�;�`/��j�yL�I	Y]�Ә�h0z�)�I�E�������x䤪�E�c�14!ݣ���n�p���(qU��9�56�t����"� A�w�������}iԢ-e�-���?2F����!^ǟ,�4U��j�l�M����^�S���V&:�V�D�����a����5H��~��v�H�LG,��>$?��,5e'�t2�N�/�m��@[����:��lk\lc�d�-��N�^����� [�<��Tv�w�g����Q��$�?�i��'J�0|����P&E������j.Y6��J�����^�J��Si�2���+� Ф�'��D|��ܹ��z���úN_ƛz���j�>A6x?��8��nxӺ���vH]� �Zv{����/�&�b���a���D-�3]#���xa��x(�3�X3`��Y����n(�$]8��;!Oֻk&G�)?yx�c=܎���?�C���wY������ag#�,��xz�M��&�QW?��%��6�J�]���w�\��(��`zu���{��y������Z�8�c����-R�Ӕ���ݔ��z����:�F�!g��!D`��&�!�(Ύ�F�#u|�; ��	�/VT	N�g��4&����Q��(ѕx�'2�3z�#ch�Q�䵼��J{
���w�mA Lg���I����J#��L�c�o���#�׾,k�Y�źq�{2�Ɂ�����z���>e��</ol�{� ��eq�t�|<��Un���T�Πz�*�ek�4��roa�mj9�\p�c]����2�W5Y�m���Dw�d���$|9g��]���/w��>�?�Ń�	]�V}�+�D���Ÿa���6���:�1Hl��'�h��@��3]c/eY�_���5��k���V$�(lA]��O/1-�����-�����b �<�����3��X5�:�:k�3ep�%5���}�ɿCn�S�;&9�ߡ��2�O��oi�6�����t����Gfp��.�[�gAa��s��������"o���_���F�<�>�gU�J�v"j����
,��d�*�R8=��k�6����g
N�^|���[�5&i�b=���z=���ƣ����X�$�	���_��Ҟ��I�~b�W�{p5�lK�ys"aruP�!?����l7&)6Ң����)"�=�7��47�~����\�����"��ގm����ZC7�ϖ�׿Nc�3�!7ߙ��e���9%U^_��ɊȄ�<ޔP�+�֟�o��S�g%I������3Z���GT(~�I}��?N�ؕ�R�?̚��栫ߨfwJ���Nt-����{�J{E1PCot&^���$��o�b1Y�n1������wx����==��X^��7O
«��9�b��6��V��}�n[z>Ps�`�Փ��l2P��J��
�J{n��@��q���ܛ�F��F�P��H���
~ .,�)�s���j1��n3�d�J1˖�*�匏m2�;b�f��V󟗺����h�������ˮ��
@�3���Y�dJ�$����t#DD��OmO�b��X�j��~�r.o#*�	giz7D\ra�������:�����������Z�F:U��ʊ���M�|�Ws���:�!w.g�Z�ۺ�
�1�)Sx���a��?h5F^ D���7�X]P��#)h������i�1^I0�$$4�dY��k�vp�>�Y�FLy��] j���W���>��=)y�q~GSL'�Gmqvt�st��"�C�����C���`	?�i6,�I��󛲪���A)C�I�>�
����eFW���i/̜=,�)�����fݬ��쾮�fP��F��b��#�^X��;=�M\������`2x�[�$���4�{#5A����������2�.I����2U=5�Ͽ����e�:� Q�ok'm=��n�_Z���pj�1 a�:U%}�Щ*�I��5�~UvD�5��|�'��G�
���OLrf���=�.����ZJP#X���b��Zyu ������{z��>	ʃ��ոG?L�G-Z�H)��i����AS�Ύ�d��C�G��dU�}�1B�|<��	N�+X#�&㉤��}K�� �\گ�_2��w��]~v��3��q��ӳ'k��yT�'[W[O�:r}7�� e�u�2y��/�.�l
@������.a}�]���Ao���n�4d�S;��*�4̝���>@pN���y`	���5r�O*����t�{y� hI��?i����$���D����n\`��=�2+��/g�^��n\aoi;~�_��Fd��^�	�G���ꄰ�p��Ə1ׁ����9r&��̺_1 Cﲢ��
&v�L(	@L.���%W�13���w>ZO���9��(DK���"7&�i@���ܿNys�fj�w ��(��g�rnd�R����8��:��������>�J ��Zh���h�Di��ӊ=T�7J�{��.�(jV�K$��!���`��������3"�.o�"~����ڤI���vlN���|�0Gz���R��:���w��00���@'�,���!g��ى�-�TI?�l�����s���O��0�:�F�����Ze���_+�q�K���WM,ڮ\�5�ׁ0:yå0���Vͳ�%��Gã��$qJ��x��]?��I� �^�_�+pt
!d�ͱH<����	�W{�3iRS�/uq���F��u���%��(SNJ
gB��-N���y+�}f}�zM�Pm�6S��n( �Ϣ���+�i*��g7�� U��d��(���/�=5� �WJ���kp5����K,I�+�׈s=?]�Ճ�z�q��qbF?���;��3)YpEk�p3B��ތMR{�:��d3�x�,?�����s�@���Z�aw�mwh=ȡ���!���V)���`Zntt-��Ώ5�fw>������o���4lm..6bBjQ��ܔa�9rt@�x�d��ۋ[wlOY3�l���5���7�
���h�Ǉ7�p�������r��?͹O]H8VO���vb����W-��L:�*�oT���0�,��W��ߘE,{5FF����<e#j���P��>�5.U-�������g����1���@�{ZMp���f\��d4٧���y>�J1/I_P�D�1z�����m�~j�H"N3�q�t>Q��ѕ��5b,Dkʄxy�ɓ���똌�#�ǡ���t��"�(�~տ:mxE�MH7��=����Qt��ѝ=͆2nD��QKɆ=�1�UKör�'��qJ���
8�Si����*t$o�s��:�~�֥N�S��4d�p�xD�A�|�}�W����W������':�E���FA	��o݅v����{~�K���z��#�(]�J��x�t��	e�P��~�B��BP��Y�9Hj7V��x6*g'���\����>�U�}��5����_���<v��סZs�ڂ�T)+L�AM�~PH��/�����u։�j��y�?��Pb�=0 �L ��G���k�������TsR�t�p��X0a'�}��4I��T�|ND<i�7��Fo��������|7�S�y��?)�$�mk��R�L��Z��)���z/S�o����8'X��G�6'�SQ2Ň�iy�ks�S��&���Ƌ�߈|�v�3��{p�x2�,Z�/s�8����b�Z�9!��\N��������:{�s���~��⹘6���2��&N�{T�Ē	��hV"�W�}���r�HV9Z�$�*��yֿ���� �Q�j��I{���z\��%H�Wx-�7�wLKV���4��8bQ�j�L�<J1rq�o��<�d�\_¥������i@�����#2���"��Jj���]a�%���ցB�Bȍ��K�E�%�/3�a��E���뎌�ж�ݻ/G�m.�yA����?� щFD%�]Z"�mda���P���"*$`<�� �;�9m|In;�1�{�5�&F�Ys�M[8��x¸���ސ�1��}z���s2ȶ)jcfQ:"�=�]~[��!��];���d������?��l��.�����*���H����a�����ݸ"����<�,��s��V�\���oO(�=¹��,)��J} q�2o�����>9�)�|BA^����cjW�xC(�æNAa_���md �_ZS�����|�j���d�|�(�=��6M��!_W�o��ۜ�a��@՞�׋�෠�bv�`�Q��_--#K���9\dt�j/U;j�Z3F���]�����o_E���A[�FQz=�&��[r.7�9�\kG
�A������:X�`��~����8�g� J qx���X�J�nb�_*0aU�m��3?_I����,s�I5ͼV�z;����^��3)�x��s�V��K� �Z��?I���.!b;���+�k�R"�w�jċ����	��I'L�)5ZT�0�F��=�Fy�����o'���������� �(SB���D�##�;T}��v~���P���̹��/�������U���&�J�^�ނ��?� �.q�Ʈ���>�)G[�ϻ����LGke���q����\�ӍSϔ#X�1�U�Xr�1�Fɱ�:`\nx_Va�b�̇��􊻲~��i�����!��(%>���o3#X��ʙ)���jז�����߄�[�wtg9U�}����.w'ؘ]����27w��(5�w�缀_7�U��O���h��a��m#���ϕ��̖qjG@��a�,����#���>���A�v�BO@L�dV�sl��º��q!��z�wI}����3l#$G,�8�{,�����o@8c3��A�?�����[�[�m�_n\�oJ�7�S�>��[�N=�!氏��iq��Z�%a�Vh�����&d�^�P�[��HF�%�f�cV��2��E�N���c��V6p/������l�a���[�/��a����������[	2�ka��k��f��;�j<s�E�}G�k�"sj�C��#��q�L7Ă���Ѱ���o��� ~QdC;L��w�f󏆍@ ���1r?r:AH�rCa�C;8�%�'�h�L�L����{*��o�@Dt�Ies���l�:�}�9�"�$h��t�NwRXZI���$�cv��ч����I�5͍��s9�B�~��m������O���I�Z&ݢ��v�U�Շm���[A	�0ha�8@���t��r�4�!6)g�L���bNyA�֝�/�s��^��ү|O�� ��L��*=�4t|��j* ���RxN*uŒ���}Q���봞*� ���v���mZ����v��ݦrM���U��f�1�����X'}��V��Eh��8Z��d��Q�Cf !���G�4��߷�`� ��R�{R=�FVv~7����|0Y��gEU���H$"ǡd�,��Cק(�74�b�듇+���>&7�IZ�MvZ��ڣ����������!�F�I'm�2Sﻡ��&�w�g�kL�I�����%X���װ �h~d�s�����H�מO�7*�a�?���YV�rw��8�����7i�s6�E �j��4���8fh)��Οz��׳s�p[����\�u�Pa;-���X	ZX�6	<�*C����H���U�	����-a+�A��H�@ta�E�n�ud ��z�=D]+�u���^<b�%��n�
\t�_ܛ�@�f����:���O�[9������-�m���su�B�TO .E:)�OIP+�G$S�����`/m-�I�r��'v͈��ڍ��� ��D]�Y�D� �Z�v��_P݀Y�cCr��g_�&�#L�8��'�>��A��oL?"gE�ť6q�N���9C����e�����ц?)���.���S�"��96f���;[vA�/�IF�����D8e-w��9���:����O~��ۋRL~g#��XO
0���i�y�RW��	�hV�ӭ
�:���{���}L����`��4�HI-ڭ�1[��օT�l�J�#�2�X�v�#��z���`B�6����D-���!Hi��ɧo�f1_r`�����U@j&M�YZ�nٳ
�'�3#
[���p��8E��bT�o��f��ƌJ����c}��O�Z�b�T��HK��E�8�N��ZA�&cu 2 ���FL6v)_GF$-�� ~D�8߿��~j���Ů>d�9����⮡8S<��3w�~=SK�	�.���Oe���X����oĽAb	H��x�J��;�N������)�ݢL��u�_d_�*x�(ĝ~�f���J�Ƚj^�N�,��Ci�o����S�#�f9UX�e<2�����`�طIe��.���x�x�<��L�iz��;�C7�g�ZN�Yo�0J�Ț�P���*Y���I�>:���ju���M����t�������|��)&�w:L1{.?����׃���J���S�_�j���il��c,�I)	��Ӝ@n'?Q�6��(�N�g��ACw�M�ly?�3wûQ�fT\�����h��T��O"y]�"��⫷�=�m�I��`�1e��m�oh�7�W��*�`���a�?��>��{Ya�6x�msSz̵V$�'�u?�;����w(�
(�hν�[s鶒D0pk>�2�j�[13�E�%1�qN�zU��Z5����U �)�Jg�K̳@�An��`�ޖ�:p~eX_Y�Q5��_�y���>kEn���&n!\�]��l���G�xU$��3*	����5��!��~U����q],B��n�釘�4�n����Jy�ދ�W��i�i�{%���J�[�,)0���Vꨇ��8�bi��8�JZj�O��&:��z��;��Y�)=΢�z8�\��f7��������\���'��I}�'�Ļ1����P`�7QL%v_�@{��{� -`N�G�0���}rϽ^4���q^9%M��]�q��ܓ�XHmPI����[�(�[�L�<���^�䮊ܓK�)�<�]-K]�߻Or%D1�')����:����;\�4���eS����`f/Zvx�B��N�����1!��B�5>���_�y��o~�\����^�.�SQ�JFT�M�#Cd�6����I�T���%N{S�A�4��C��rX+"@M���q�{'s�Dw_,n*`�?��-X���8�ͻ0�e��ۈ�ܖŉS��Kqq�8�j��l���
�à<�F�ԙ���pE�NP��I\�Waקt]��4��+��R��I4�勆.�����hN�8�~����Ĺ��I�4l���x���Z|��/��@#�W�q+�&U+t\�Y���� n�K5��jՐ�6gS��0�N�]"Џ�hգ��!vU;����i�*�0�9�c-�	��\�S�W��%�p�?�z,�8��Ҭ����W+���P<I��ȕ 4�,d�_�5 k��-Ε�i�@0��	"�OT�*[Si䜁G���j�	���%�AE-��Em���E��"O?hB��Q�.�虜v�` h�)~�ôፂ+�#
T�h�`eڭ��CV�h��C��,��,�����׬R���7d��%��?��q-�>�u����$��<)��G�;�8���H:�c/>,�+�減F�KUf�D�3�\q�_5�p,��/̕KL��zQ":�$�9�
ޖ��v��� ��tP��Pc���6	 ��>�k��C��2nj���N��T���B�=R,ع��r�*mRyk���q������¡�~�D�pt������c��f�k�Ϙr�/f�ݼ1qiH���6Y�sR��p�Y��R��i�k�[�֦��x)jS���"��A��DD�*�F(&ob\mW��ơ��e�3��"GkM�m�ŸMc���ڎA�Xn�˜�b�T����I��CF$$��9�q=O;�ݘ�I�4q�\����*�7v�Lb����)�N㵅$o ����� �NU�'��D���3Ȇf%
��Z4<��FȣL�n�R�J�mG��O�:��h]�5�y����ۦ�Ӡ�����^j?R9��ۍ@Gɦ�U[N@��Z��W��P\qY����O)~�FnJS��R��P��^�LƄBC�l��GSN��9b�(��=t��DJ$\7ǥ��y�����7���Uva0�vc��Ѻ�W�ō|���@2���Xe�h2�:ǄBbd��%ic�tZWZ��J
���ƛ�~mM)K^<��_N�jζ�_gn?y�,�$�.��dW/^�1�݉ީB��l�;���k�`٪
+���>9����O"�G�0&�5I���Gm�t4���l��"��v4��_����'T8���":�v�C��O�B�R���L6o�c��r�z�ދ��S,��'�}Wҏ'��Q�g��{I���b��t �k|�u�AS��|�_݆��_��6x�g���$����[_�kG[���i��Gw�1��\��J��K�<��*�S������R�N����z�Q��)LE���(T��~�$����G�
K�lN8����=_���|�"���ϬW���9E���2���|4Ԭ�9��ؙ~�OK�*K��F�B�D�("���T�iI#��?U�	�ԛ��w���̽]_��t`�x��^c`I�g��IK)E�L���
qA�)���]��\-�ϕ��g�Z։�\r�PM��Y7�Y�C,B���� 9	:�dϦ����9b��z��D��B2�_ўK�ܥ���D��	9�]��|h`/�}�{����T�={�9-<���%����X̽��1����|�ʅ���y޽ir�.� �цh�=�+�ɲ��^%@E���r���a�zs�wT�����͖f�;����}��c���XFt(F;p�$'`������Q���Nbt��#���Z��ױ�􎀝�\��Tk���}��'U�c	:G0W1��Z��W_ �QCU���S��E��o�#*Tæ��9�ϫv���R�ߛ�?�.����
Xǒ����-N�Q����P����\�	�r�`H�:T�v��R��'%F�iX��⽿����0}�ӗkH�#�$����4��?����͉�CF��;F];�~'��_�Zo)NG��i4]��]�ݿK��T����c� )E@��Dc�o��-�,ؕOIH" �~�;���� �7��v����h�{H?|�������6	�6�6cR$���*6D­H�ѐnŒnoBf+�2���'�&�s:Უ�%/v�}k��?�d�n�AD�O�n��̻	W:,���kY�>��k��Щʕ"�Nt�Mf���t�,�B�����0�_��k����%Xw=�o
��ί�:F�iHhTjIY�j�P�V��D�7�����}��i7��$	��A����Q}:�ɘ�Ǆ~)��dDkv�0a�?VĨ��"c
�;Q����֍��hːq��"q�:�f������m�]��(�븤�F���u��e|zx����Ӑ��;8��7�i~#Ɇ`��A��E���*Ro"���2]l�6�u��q��L�_`Σ��>��*n/,}���(Esp���w篾Ҧ�������)08�ײ������[o�b8�4^Z,�a��lP��	 ��\"�×�ĥM�hZm����,A۰mT�����4�`���E)�q�!Nr��F��0;�ٿ~}0p�8��?M�\\��X�DW��>����W�JN��*CQ��w���&k��u�`�B�L�{�����Z5���k��R��%�ũka�(�@p��A8^�%f���B�G�Q�����9��-i������>!7%j{AG�S1B�b���&��� ���|�<�]&+�7����}EF��GI�G�z�M�����V'dj�Xi�,�C�޵�˿��ތ�;߻��z	B9d:�Z!G�/��]-�\��&�xZ��F�a�H�_m2'81x��
���V�חJmp��5lI��T��\>�R}��9�c���YF���K%o��}��f)sR�u,ϒ�I9��O������ �2�8w�ܺ���~�v�`N�x�̩��^��Ǜ��|��7U��c{���O��4(-M����t����!�Q��,ȓlɞ6��qTe2Sbo65d��xC��Z�˱]K�+x��P�m�"�zF�����B+��[��k��
W�SBc��*�"�9M(M��X,#F�n *%5J� �Z :�}��7���B�UȲ�*X2%β]��b�� h���<����]3�@{˦��G��<U�&�h���p
�9c�{ڔ_����2�l6�%\EQ��3�D�J��G!����S��b��D�/ �7��3~���o��ܒ~��Ö�W�f���Ty�1� �0��B�9��R�ϔn� �sY�r�mB����gՐ ;�㍖�ΎJ����Ű���p��3��oķ��l��שk�m�J����Gof��y�l�a��מ��톖 Ŀ������g����ҷQ��&�����-�귋��+Q�gD@j`������M��<U���S+������Fj[{���G�5�o�%��ۿK�*C�$�)�Y��#V'F��A�Y ���F�%|����47)rq����j�E�\<�@V����Uh�ށ��V��Q��O��V�]��ɵ~��ܤ��3"t	��٠>׹.�qJL������|�}-����a^5��M꡵�����Ӣ��u���� /�t��'߆���Vd�zX�Aa���B����(v��=�tkuق���?�p�;���imWN�y�4(,\j�'���f�f����c�L�ɂ7�
^X�^�4�`�Avp��DF����헁���7�� ���1�>(\�ݹa�r=q���v ~3��w�&��R?K��8m\���V~c���z?��s��='
��M�_�6�;��R=��l���Oq�;�eͿߕҠ��	08��q	aR2��e�f���G�"Z�ӂ=���yfO�����%��)Ac������ʮ�������, ��9�r��I %ՠ&�O�3���Ј��'"�hco��i\�4��G�z�ZN�ݯ'(���;^�1|+�`���%����b!��Fj�SL�;���*����	�����7SNI�G�]�����bLm�IԖ<��S�S��J�ޑ����ם���mf�2�eCGA5}����g�Tk��ױ���ۻL(��*����[t[-좬�R3�:HCE8�[k��"T��2r��u{��ć��)��q�3���B]�s[����x��-���M�o�p�HH�n�o�s��ki]���՝:�x����U�谥z���%�K1o|�u}@��t��/��-�,5�A�Gѧۖ4�C����
tW�N��9�јA fo��C����:rqkNe�g���o^(1���D�cˤ�W�;�.gJ�"c�q�G�h(\n�B�Vo�.Jپ��G�]kCv�B�Ă�H�'!pGJ��d�����z\�QpK��JНᤙ��Jug�:������c�XI�UӰ	�[���e,0��!<45 �Nq���1����,����6� �"�J��V�IX��Q���)�G�ֶzz|��*:�� �aɀ�:���p/�'�I��j�$���t6U"����p"�G=cl3��܏�>\�!�n��w�o&=#ylG�n���Xw�%@(�PX�K�d_S��7ίv2ʿ���%�Hq� ���s�zɿ���9o��_�#%z\%I>W��ZF(����j�=m�K9+bM�F���,�}WhƎ(W��% x�Y��0�)���$�z����_�-��_������c�w��l-�Id���zp�n�'��k `��x�@�ߘ0��(B~i��(�j��WȔkN�4��"`ɢ!B� $i��Ì;@�����!\�|g���b��U��.O��u��+���N�Ԡ���|�u
�y���M4>M�ʆ�d�v�~�G���`h��H��p<�t?�	J�N,Bz=6��W��TqH�`~|��@�FWa�w�OS�D�	��4�4f0i�-+�f�\���RӲ])Q+�k�`�+	��>7��Z��X}�i1���˧�DbS�ʛ���_��W�(N�S�߱���%-�Q�d�ŪW�:�Zhg	������7֟��@�
�Yp~�DЕjP�׬XZ��>�z�f�zW��E`��Ί���y�����::t���p0Ư=DpH���%:��}�s���9Avh���L�a+��ٮ6n7WC� 3%��~E.�t2��\��2�� ׺G�ّA��4�����.�c�g������n!���]3N-�<W�~~&(����p��2(�0�գ~;خ5Y*�j7�ok0�6�����$�XJ� 2�y�Ibj�n�H�r�N	aO!���QV���=�Hr�t^�Qu�:�M���ӧ$�HZ��{N�]n�x	��"^xC�|��+��O�z]\}�	����?��OS`d�x:?�����d7Ͳ�,��]97E��n���C��C��:wcF9�u�hi��z؋*YK:hi1f%��ز�-��R��h*{iW"A{n��豚����xo���sRSק���5���rI��H�
�ƕ�[�zu]�W�c�\�J�/B��%�q��[�B�̗��z�X,,͛�*����ii�8����Ģ^��j�q��B.�`�1��!�۴%RT��Ê��2 ��~��KC�#��\��I<����Y���E?y��[	uX�T�.�?�3�Q����Ǆ����q9I%��5�f^�όS���M��DQ�]_T�iS��P�̷��j���WsM�5
��4�u��8󇘽�]����*iC�.��=��k.ب���Iy���:�ߠ��ݡQ�y���c���%
O5b�\�׀��/�jۍ�%�y�ߩ�a��i���S�]���Q�<@b�LC���x��I9��|�:�a~ʰ��;u�s����R`]^���PSJ�x@�������m��s�O$
+8��A��4�`��@���ʙ��ظK�s�5�Rn$�n����h~�kdУ����{��~�!3%�2!�o&��FV_ns Z������!���c����'M���� �Oh�~n,�a;_g�Z��r��Gp��oA��%#��� �~��Z����&K�;��֮쵑 S��]�y�uc��i�ӈ|�;m����j*T�z�U�2���<-H����im	1�:�g�"1Yr)Ӏ��1�-2�_)� �-E�U!O7zY.^w�/)K<����Y�]ٌ.M�F.� v��u�ѓ�[7�]�3��kɓ��u�+
c���/kq6��
����Z��;-%@�.��	Q�ֹ۠W_�!Zd�l?F;i�ƹy�U���Nb���2�_+7��}g�fp�����+p���){�f��:�Z���eX�]��|!7�(�����+�+lC�&5�y�Y0|G�X)v���v �]N��៱�(����~ƃ�Qf�A���2��)A��,��Ja��^��7i��	�)-�?9`v��'�7띾���RŊ���c�����Ԑ��}@������pj�����{x1�Y0�D1�y��):ç��d��q_Dfh�d+�^Yh�/g��A�u!2�r�M��y�V#���>�0��m����ѽ����-&�u���*��x��I�jB(Xܚ����n;dQp��sH�&����#(U��v\�4	���m���1~0��v��hw��XhN��ş��"/�_r��u/�Ē�3��b��EgM�a��dM�2,���i��X�G^B���ޝ0!Ԏ�Gz~�z�'�M�Q�D�}2�J�#FUf�80��?�xa$�~�~V).@ ��dJ����<ٶ�L�������h�{]������s��R7��쭃��pU>�ĭ�>b��1pT#^Z�EYZ9�O��y��>�{r��<s)A�q�%/M�X?B��!��3>�&�Ls���h�?�H�Cؽ���%��e_��-��!����A�7� 3�-�]Hoo���BkQ�1���S_=�(�5���g��K�2�K��ՂQ�x\��.f>��+m����wG,�/���Ŕ7_V��31�3�Ũ�*��W�5l�{�N����b����i���H%���j�e%>zز+|�f"��w��r)T��p��'2%h�74(f�_��n����J�ѕٞ<{��"��I�f���E.��fp���g������t�^J����6�a+{t|�8h_[��S.}�����7EKV�p��絯N!,Ӻ�wñ�ݕ�U�˪��3�����}��O�^��@�*L?�~�j7�����(�:���%�Y�L|vf�F.����Q�eƪ?�=+����TP�`S�\=�P���J|'��mN� ��[A.A�X�(����;��[<X������x�\���*Au��"� 4�~�16	yE�#'��:�7#�O�C��W?x����<+��f;�����S�jif�/�
��S�z	׸8ÿ�֏d�c"hɞ�ڢ��+
.��.~��NR7�z���Z�}8%bɸ����u�s��(��Ά����ej��t��/ ��ҫ��2^�(�b��^�q-�tc�P�!:O��r�@�zG��ؙ��3�~䃒zp��:&)@�[��:�LS����{����TȇEe,�Ą�w��)}������/��͟~���������}�:S��J}���$*��F�J��?d�T�]�-LKq���S�]
�P�ݡ8���-�Z�]����Z܃��~���ެ�E��9{�����<	���`� u]v5Jh���m���"Y�Y�ra��(:��d�$Ƚ	�5�7�D��M/6�x���2@���zcj���K����G)�/Ǎ�*y��#.rȲ~��S�;ώ�9��ʼ���K��@1.sD���3-(��o��`c�DА{�?d��ۯ��	"��6��-�"
;8��=Q}�^'$&�HV)���eF]d�>��������Zm�*��B��~��F�Y�9a{~��Z�������P y��8���(��MPg�D�NC>j�80�.�@cQ�^���'����4�Z,�
*�kѥ�օ���9>_�\������m*����j ��m�c��#Ǐ4w��?����N˴4q��o�\�E�Wll�jG?	7�w�"Y�w��Qَ�I�[�f\f�Ϟi�=��g�u㐈���{���f65�~�	;<�V���w��������d[&Z�ߐƔQU��4#�(-��C���4�$��j��B�Y�8���4�� s�����+o��~��W:?t�������i>�&�c�/����e?Wϴ��~=�ǝ��NbS�G����g,�~1�v���H�ڡ� �vMG`�[)����q�+��7�����Nk:��j0�5����e�G\��Z�h,ߒt��]�(F��"�y��q��V��L' �!��d�.�����3K��� 3� k�%ȣ����ꉛ<��Ȓ�⊝��>�IRO�r�<g#c�-?��P4���Y���M�9������]��l\�Ÿ,��V�x�zHL�E^�~+����B,b#䌃&�1��Y�b�E�w��y������rLxU�%k�O��*�뒄�'�MfJ��h��Or|����Y��m	^��Y����Lu8��)q3}\ߦ[V���Þ�<����a�W�5�f�sVZ�$��ݹ�CZ��w(���W1������x� ��7AT�rlT����0�q��D�P"|u�~
P�ʻ@�6�q��o��J�H��p���k�C�v���5 ���s⢤@��)\��u-���O��H�[��SϠ�Zr�!u���xH��AV	^G����!j�ԃ(!C��l����w���:��o�y s�u}���\Hһ� Qi����sѵ��y�3���)^�g�o�/�B��4�W]�����$@N[�DsW�"�
CZ��r� $)��L�<R܊���~fƴ��AK��������:��[�}��`~�4����/s��-�����40y���W������2|���Uꬌ�G�:H]$G9�Y	���W(6����59�������G����j r��a�9&�_��W�-p���-	 ���X��[����7�/QZ�����%}F�����UW���Ţ�@uڤ��v�I�^q����V-�Br����F^`l8?����(e^4��d꙼���[�h�ɡ\�����y��]"|W+����c]�8�O[J��K_�梿��߬�?�BS����mty�AR���!�d���p*���0��-I�o��uJ!�0g��n�?-
Oz 9V}zy�CD`'��ܹ�@D/�����&�u������Q�]
Z�8��#%���ܬC�VI
$n�`U�X6�M���Qx��R�ʗL�d�̻��+=�񰳤?5��K=%����IR�Q
� *W�U�>%Ѣ!��%w�)�-З2O����]00ϕ�����P8��F?�EDEX��\�>S�+���wq�^���{�pё���٠��'�S���IĞJ��ZȜ_ix������b`���Jv>:R����P�axUJ��Gc��H�4�hiE/W�������C�[�25=A9G�^BF��/~GC���c��l[����r�|`H|y�c��h���T�ʹK�:8cM�;���5)��q%�9���3b��y��y����O�2�<�6�������=�{i���f�Thm!�9ou#�Kv�E;XQ�K�aEw�nS�K��Bv7��[��6o��.{	]L���<�|Ѳ�[��)D����뷣�	��Mn���n%���*���~%gQ��},'rƶ4S.���Y�͞�[񳙗hHV+Dh�ЫΡ���x'��(��.�'��Or��a@�[�NRiI�aJ��tȂʓ����;A�<��^+�1��A�[� ���H��#D�|��%�/Cl���.�� 
�n�5���{+!�����&mA�~����
��M���a��A�o-<۹J-�
�YҖ�� ��zg%�TAp�����s'x�R<h�5l��N�3H�L���Td�R�4���˛�J��o���`��V�;E�;^�b�������ؑ���-�/"�ɱ<[��v����I�8� 1�[�&a���xS���M�ŉ��OG��TiE?!1���x���0���E�j���nR�RC35J��� �Ț�-d��;�>z���~S��c�}r�iu>a?����vo�&j��~��AÖ<W��s�_4�S��6�q���n�L��H�^V�jq�#?ycW���MƵ6T"�:,N<�^~]�e���z�J�����A[ ��لqozt�W{�_@\ ��i�^Юn��N���dwoA�����8K����&d5�Jz�oLk��F�HS�zr4����4�m��4)��Z�}r��'ѱ����_'T�^�YO�ep6��r��{��Q����|�H�NE�P��q,5]|�娂��I��8<��x�X��Q�%c=���� ���h�le=�n�S���iEp�y��p�?G�yZ���[63�vy��M;�`�z��V�d�S$Ym^�W�.����AZb�;�h�k��Ԡ��M��O���L�n	��#\ӭg�t��$�����97��Pxę"�o��v�+?� Ь*1���tYZ^���
�]�����;u�Ǯ��`aAЇ��kz��.�+2���ӄ��޻
�G�9͠��8���7��|�F���QO�0�t=��ס4��.���x����]W
�%1<��F���=��ϋ�y���5�7������+ZS=���h�X�F�<<�%��f���[w-������K�Q(���e�NK���h�u�O��G�Ztg�-R�,R�Ń���ɴ�ʜ��Jw���bsީ*цN0��/K�kN}�
��l>�Sgm�т.u�`��5�W�BM7���Փ�|n�,YZ�&��8:r�qpbIX��V��F���6��O�z;+}"��ž���	ͅ���LћV��@wu:�$�4���[��}�f�D�w��ꆖ���zF'v=7� ��e^��)A�uX�v]��Y9�ڼ�� -�t������sK竬m�aq5놪V� 6� �2b��RaI:��_o_�jW.��1�A���U�Q8�*�P��Gw���[�����w��<����)ƉWJ0k�ׯ���{IB�g� ��hgQDY�13�A����uʛ�X�e�O���W�����8�F��c(���h/g5��e����3e�H@�Tcҧ���ע�����`�JV"V��E���9���>X�Y�4S}�A�0�_h���1�)��t�[:�o�K�)�bp��&2�g|n\�VW��b���B'�KX[{�Y?t��`��zǵm���|<��Ӓ5�r/#��6Я�e�!xÕ���x�	cFef�?_�y�u��?��O�l�#�-e��� s�Џ�v��=ז�Q����T���]���H]�,�Ǯ~?���>d��
J��\�o~��hp'L
W�
��[ ��v�ť�"S��\ -�9��� �N�^ςRn��3Y��`�02�`ba���,�1��V�����к�7m%ɹ�Ի�w߱��xH�����S����"_!�)�z%�5�#���Y��l�=�3�nz�jL� D�}\X�ˌ{Y�D�+����h��8Fy��������'��լ�g4Xs�������c2�����b����z�V��@�T�?�LW�´���v/y<���G�y�=\����\�,VC���J*\���[r碫�O��"���^B��t��D"��9Ok���ɟ%V�{�*?|}�P��;���;v'���
��T��_p0GvI�z�8N]d4����뎶�J=��66j<���:.�]�]�5�8#F"M.>� *�,L�7�;FԸ��=�&$���&a�9:�;��h&��%]��B����$$����jv\��F�J'��"Ύ�����%��k�uo�)���c�g9��p׀�S�z8e�Q4l�z��>�|���pl���B�� g��i�K�Z�%�у���y�zj0����;��͇�F��u|� -�΢m�c�ݬc�Aү��5-!������Y��lӚ}��{�aE�BC��ۯ�`Z�g�ou�+�=g9v��<V�l�Eg\�ܟ������g�q��X%=P.���_����o�`�+��Ɩ�%�ሥ��F6������V[��l��nI.T��2R��U�^�eObZ���N�|�5��e���i�m��W�g�W0�*�¥x���֎o�����NY���ك/�`@>c�uc��-x|Z�F{TX��VeS�.p.���R��}0��H�L�	���n ǌ�x`�ap����%�=x]�ٕ L�x:}�+a��4m5ˢ�ÓV�=��P���
�bS�]
X�DnU�0���9�r�L����Fol<�d�[<J!��}�I��0�����g��i�{}����ϵ� �4s ��~#x�|B��v�}�����8��#�k��	�%�Fy�j�-R��T��&�KZ�t��0�����P"��kTi0ź�Ǉ8��R1�� @$�[�n8����_�C��A5g��9d�X�z�E�P�!!�{3&&p;G���.q��̑��,��q���r��R�8{b��!DȍH�i���n���#�D��L#������k)�ȵ�����#Yt�6߈�<tH4�K�ƥY��cv����vy27���\�B�&G�N$���i�/-���u��{��U�~]���U�YYl[�t��Z��|n��2u��n.�p=�6u�tR��b�ݐ��~9���B�XB���l˕
��c�4�8~;gT�S�ծ��V﷐����7�녵��F?�Bc�2=N�s��&kv6(�Nɴ���>q}����Jf�:~R�D��IX*�����/��j������f"�J8p2�\q�l��)��D��;HÌ��@��9�f�0�;`֨��o�ʁ�~"c]|��\[9��U�B��v�GǪw��?
���3�or�!L}��X"᷺�
��ȑ�ᑽ�x\��N.����fU�(;�u�M�5��ɱ"O� ��� �nHW�5d		�M�)ROC��H�k=�N]l� *���!�f�+��P>Z����RyGj۳ż��GL)'���=�{т?�ڜf�{霛y#۟�Ei�m�Y��-x���	��K���l���I;���F�;6�����������Sw[���E�X+��I_�{
״����e�:
_gAa�ʴ����^�ŅC
��;�7������� �?@�r!�]?}Ü���Z��{�sӖYJ$����R����l%���6�T�o��������#��n2���C��X�U���w�A�@�k`ےі�3�����8�:[�~��5#���j1�@�y2����f��<:���:!���K��=�L��t�$��_�;���S��\�w
��mh�h'���k@K�
y猲k{��-R�0�L#���
�RT��إ����Zx1���W���0�s��{��`h��G�V���� �����K#F����}�d"���Ƿ��+�#5�jp�FO��ij�D?#�I�TZjDmӏ雛љ7.OsR�2��36ZN;���������4|���Ѓ�T	e��`a�OX%�%{!��H���ݘ�VP 4�C4*b
pvv��!�6��HJ�k�ކ۷�a������.n��<�LMp b"���xI�4jn5|	g�)����W;û�� ��nf���Z�JZ=��� ��Ot��C	#�Y +� ˨:WA�\ �)1��ZЊL�;�[P��/"���,ū묽��Yo�F2�?��6���ـlސ��t��M�:�'���y�'Q����z�X�]׶���� ��*�����S�KN� 7�'u�{H�֪<��*sXf!mw�M��{�������[]o���ĩ�d�5o#�!��4W7,�s=~c����a��$�2[�]�~�Gn$Y�wi[o��T<�ʵ2'��h��ZW����\���.�XW��+RG�Sʾj��Y��'`����e
MS	���Q�'�i��S�Ê�X�L#�yg��(n,O�V��(X�X��F�M����JRd[�E�i�V�i<�>�8�Cz^g���ml��ث�jm�Omtp���
=�=��h��C�m�鐔�C?�]`�> $e� ��*��x��Ar�W�j*�."=�k��Gg�#U��
a��Rn������YH��M��2�m�|����E�Ғ�7�V�ңL�@�}���O� ��q+�ΣUݯ�L¦��{[�}��U�n���}�Z�s�l�t�x�yb"{.쬵�Sʋ�]��I���0
��#�����̡�q�<!F5��8����AH�֞�ۤ,ިiX��Qy�v�m6��̀:#�l��L����$��q�9��
�ء��EZQx�<c�L�g��=D����|�l�3�R��H&,�vP��U�#ױxU��݅�9�%� �f5P��p�B�\b�>�@�cɩ�X;<��w*b�����,��P�_�D�hU^4�I�y��F۱ǣ�='�%��Z�m��K������ÝЊ�C�ԟK�Y�<����艴 ��Ⱦs��D�W�d	�#����Ǿ
ܫ)Xs=�8����J��9*8��M�D��DB�*Q��f���?�˜A�eg~�4~�Rӯ� ��b��������]����o�g ���P����L�kX)�Bs��ҖM�@�o�=�h*�x��Bce�ύ�j�-ݿ���e��LU���ڢ;��������v@�cLܜ��v�S=�������f3����:m�{ߨ^ƣ�0\3�dZ��<\t�v���p/�"��P&ɘHH�s$Ij��5��9Ue(C��kM ��paVA�g�)�����w�و�+R>Mfl���NHO����v	I�n�J���+z9������~�����3�%��,�O֚��ñ���g��L�>��]5;�`җoJ����h��ҩ�Vk��D�L�P7�{ϋ�i�n���t�P��ί��?�+�������h߳'G�V)}���?���'-JW���yDR�7�ɦU��˰dbd�����#�8?�-�}.3�y3�m��d�s!�~�6!�{ϼ<*���H�r폆{���P�~��3����"����H��yՎ=}Լ� O���YB�����ϸ�&�g�(\�����6?O&�apMM�*|�1_.>(h4~��0@2r��l��h� ���ǹ��^M��`�a�ڜUv����{]H��(ה"�:w̲b��~�уmD��&�]�/���_�c��{?����:p�嫻`��~�t��SCv�"Ay��n�CA�q	c��K�ʍ�w�������B-�sI�qij��!�AZY��ݼj��܍<���XL�}4�i��G�\�F*ٚ�r��)�Еv�HW��t�(Yiw7�]����V�l^ʼ�kh����sN.
��d�u;��:����a�_M��mH���w��I)�����Yx�#��!��x!��������Oc֣{���E<��F/��^f��т��nU<iKyZF�w,�.ey_D��<�<u�0��o���b���s��Q�;���j^D�v��/�78)`�� ��h�ŏ�܍5��}4mq�TFg����1lfI52��]���J<�]O�h�X�B=�5ʪEx���<c��Y��;�6O&<����-��d��P���[c��:Yͽ�b$�z ��'�&��z�
q�����֭/	�78x�p��5*H8;4yX!���H�|X�}�cg��&g=
T7�1;�)>ݰT�\�I1��hZ Hh:ހ��a�m�l�8K#�p�x��:���C�Uy�J�� ��`���O�ΣfF�E7��NᛦW�
�~v7Q��G�LM��B��}{���U���2z�u� ?`��Og���gp��M��ώ��Eg*u0����a��(���\�u�	���	x#v�;g.:&�����a�03"���BX�����S$�F��k������-�cF�N�C��5Doy=?}������RRi��Y�Z�u� 	B��� םa@�Ml�n�LxJ�1m9�^TQp<ޢ+��jcm���`1A=��?�y�VQ��|�3��|^`��}�Td���:]&0���W�
�h C��ib�9F��X�7�¿�_(�F�=۰�[R��L;�ڼ�nC�wo�#��#��ݴ6��f���QN��M��zr��V�:��)��!�ÍD-������$�6�/�$�K<�l���:��[,���nz�~��i��Er�R�b�z��I�sFٮ�54��2���8�#�[��K	��M��%��=�b|�z�-�J�1Q��F��=U[v�8��9�zY�����t��V`/�^�W��7��ӏ&����k7i��>�T�?�I3k�^�p*���+(�$=g��9Y���c=��~�[z�U��x�d�I2��B�~��y��匓M�GFA`d.��t��:�
�s��k���v��gA�Iw��M����z��w�ܴ������'>W���5�kA�NĲ�{؈�v��c����]Gm�BE���.	�B��,Q}��ܽT>*r�BǨ!��7��u��{���'s�A<Gn�״�R��D���_L�G��y�;	eD��)��uB+1
����CcR����O�PK�7L�k��Db��� ���  H �	��ms�i+B�Sܺ�G4�Z��^Kh��D{����G�Ʋ�ݙ�ŭ3:���Y�'��Ì�`zA �>rsR,�[��������U�C�͡��i���M⟓�Ք4��X�f┻��?l�R`4�C�l12��"4�g�� �H�Yz|��k��zۮV���U�B�/�-��jPa�Ң��:�4�@��?�3C1�}�ԛlnT�L���$�|�c�ѱ��Ħ��(��
ۭVa�ed>K�O�}|���]N.n�π���^�u��m'_�@æv$�~6K�W�|؄�k���=zm�0��e�5�I)z��>]�B<u�5>g%��k.O׫��<��h\�Vn[$�\��ӣ3zO��O9�\H^n<0�����
Z�	Z�d�����o��-�py���7'q����'�O$K�RS�對�Z�0zP����Ąx͗�����5v����t���f}9F��p�t�
�)d�s���t��tqW:�g��pl����B����e|LMH��N9�1���Xd�B�l���x�Y��1G\�� �꿚��R��&���G\~}���P�\�3�@%���l�����p0�t���hZǗ�����G8b��C<�0>0�'�k��Y��'�CU�Qa��O>��|����o���M=l:^���g|M�!*��6�9��OI�%������
�?cqȐ(������o���d]o<�h��V���6=�X�1�>6^��&�{������i�*	��T�`]������������}̞���eR-�@�Y&C�{v�+�_�\#��P�Xji��m��W�V+s�6r^sW.:�kN�<��z6h�o��D�}�X�W�,�ƥfz�]�;�t)��rI�!��DI�}y�m���H(�W�{85���M�kw����=[�������w�t�dI�517��*T�!��&E��O
�Oi�d�d��������D1_ƙ���w�~"�@�y<_�w�	lw��C�yko��ޑ����o3��>��G�G=�Q�q������i�V-|�Y��Y�(ՠ�QE�8�L��f��j��zy�5������'|�)����Mv�~�C�x˒#6Z���A(�ۿ���nYs:Ʒ?�<��=�������?�::�@��Q����D�r(ֆ3b	�H�m����-i��yտ��z��ҳ�[C�f˚�3h�I� ���)��@b\P�1&�$�V��{�v���S��g/·���'��@�C/����������n&�Z�Ów.=��>g��@�R��E]��n�(#N�=' �𦇪-�3�U���ߗ��E��@w|���2���y
��|�qwF�hݨN�����OR۹L��o?J3�h���r����}�j�z��QW�}bF20������/��jI}m;�s ���z��8�����񷕞r�|�#3�0�X���@A��`I�kQL�-�����q��FPqZ~"JUGm��R���x��G��������T�=U��o�E�~�]{%�c0�C2K�7�C��=���;r����[��p��_Р�F�ƒ�o���6�-�N߼������N	�%����5���bBˤ-��.�m��_�RM��1����r[ۆ-���RJ�U�*f;�_,��7ͼr��� �i�nON��t;�Ϙ��f+��3���|�_�2����D��D��
K�� Ōg�Mѩ/�ZOs��|+����cy[H��|�����'+g�:{��!�{���w��̧�O�ZV�8%o�q�B8� �D?����l�(�K"œ���(d� �s��4zT��v�b��CPm��9.�:��ox0��u�F�+��/��׺�<�e��g�'��7�OE�	�u�>�.��\Ԝ�<[�c�ƺ�P���0N����7�2�e6{�m�����@�� ���2��t�+�\S6���E�����g�C�9�\���!ӭ��.R�Q�Ё�{�\��C���$��y��b$���>�y
C% �̩��8�g/{��+޽��m�a¯j��{�O����2D�21�p��|R�j�C������V�\
�ot�98��e �]�puC��#s�`���
*�l����r>D��͆ �f��P�\��&�k��&��]zb(�wzXp����Aْ�,���$#�*Z��B����7]t�Ǹj>Z��[�sJa���-��9Gp���uWC9�+��R¯^
5NJ@��7o�A	�n`�e����֣y�N�<��=�����菓�8#GB;��]k��G��̟�9���87R����'��Cn�����Yʀ@�X~.b����q_�}Jk���QKs!gG���2�b���D�����	���.�h�xo��s���]�u�@k�h��t�B��ѩP���WX;Q��Ȓ)I���9#yɴ�mka�us�d�ϧ���`�2-�K�'��N����T<ש����H��M�:�?&�z��|��ם�4�S��d~���d��L�I�]���V�U�9?�Cuk�Qk���b�c�%��o6W�J�o�3yC�^��Wn��^�̘�Cfq����5�}&ts�S�}��Q��9~�|��Єt�@G�ĥ��5O���,~	CUs1[9�������C�/��?���GݍV�������GK*`5]�#=_˺M���kY�\����tN���	�m
�\�x,V(����~�}#j�t�q�@C[nM"NoG���֔&q(�q�ܹ
����"�_����۸%��wfvT�[���űl�/.>���Y �u�m�����뇃�G���p7�Oe����AG�z�w�s�j�w�5?�y:� �;E]���Q����S������E�W������}]#G�ͦc%���rw�h�����a�3�S��E�[,%mݟ��,|�fE�k�h	۵;	�z���S/�W���1���s���Q)�|,5y� �E������я<[j�p˯��oOܶ���q���EDAX7N�ن�]�tuR�qi%\R8�np{W�b�Z�"�oYA�D��,J���+��;�)�F>+�&��_��s�H�w��.�N�A�}��mF���������[�UX��D���w\g�q����L���ܜ���d␳�Z��Ā	c�qϟ���o�U}������x9w���dl�h�U��z096����/+b��������4�~�)�T9:�eOSe�Pz��v:��m*@`�����(���� /*�7�I�[)��D��C"��l���j�^�����S뭐V��3���<X�xO�I�I ���k�E�֡S{���6��;�*8�?PG�>>-°��1O8�s�Ō�lG�w�XJ�.���$�I����m`US�E��M��i�@u�o]j̰>-�'����&mMu�?�VF*�գ���黺�o�s��Z����,G��2k��B�t�t����V���؝:y;���:�nd��P	%��Q������V��~;&� ���FI�����!�` �Be�[Ԕ�h�U��q��6PeF��!L���A��S7gf�H��x���?�j܈���]����_�/#wWz�t=�5]82��>n��?���L7L�ֱT�(O�]1�
/�ᦳ	��x��Y�!yV�Y/
p1�[fs����>}���s\���g���	���p/�_���*��F�AI��D��d5DְJR����:�8�Mw���/����*���e8��4��]:�1T�(�ʿ ��1�Qȡgp+F[�"��,��b� �+(�8����#ݶ�_-�e�'�j��qRE2|k��?��F���<*�j�M7�+�����z/�����NO=
1�?Y��qf�H�2��i�lRca?')�t76�\�ls���Oυ��Ѯ��4���͏)T�..z�H����W��".k����|�RSdr+ǘ���sQ�$G�B}Xtr8[#+���!Q1վc�bbk��ʫ���ӅsNg��������.�2���w�*�K�(�*�W���_��d�RF��by̵S���VX�Ge~�<|�]�xe��E2�C{�'s2�#��@���S���ja���ԑÉ��J;�?���w��g'χ�Y�ֲ���g�c�f�0Q�3�������E�V���
,q	�% ��H\;MK�:����N�|�n��D۱��;̡A[\pbU��c�]	��z����R���ޓײ�"&��K�=��g���I�4.F���$D'�</m8�k�t�i��9?��p���P6��6���%����D���f����z��֌�Q��]"Έ�ݵ/���&[���ߚF�nG5���sd�ь��z`���՜0m�E�֍?ht(Tj|�b�6�d�y������2���G݊����d��L2���?1:�#�S�k�df��m2ۛ,�#C��>�f���[i�fO�m���@�>����>���B�{�b����U}߅�E>@[.�B�Ib3��:q��'��a�fb~xjV�Z��\�T<�ΐ��a��Zl?�2O�����'�-��r��{2���>T��>|�?�¹�q6}���|. Q��P.Hn&��!�輵��f/ަ&�2P�����k��ri�ގW�D���0s+sbSr�ϔLG�O�J�8A�Q2K ~gɡr�Vۼ�	��t)�����A�j$~��#w E���{�aX;�QZ�Aڀj"��?I����Q
�Ԍ�^�hi�;��Q?M���ͪ�^iڎ�6꾝�ѤΪ4r���ic�HY�:����������x&��\�ˠ��{��z.'d��묛�f��lZ6rQ���^:�(0�O�H�	Ӻ񷽦A�$�Ug�	���KWm��`vx���z�	7x�N�}besƘ���:��M�2T�0����k�7SB���e��]$�ƶG�Ƞ2M�dR7p۟�	�G�u|TK��e�ں]�L�2�
HNSp�ۈ���+���]�U���4�tm\�DO�E�;{��@3�B<��U[7�G١�E��nTj�Tk:[g�v0Q10�jO��t΁ɼ�V82�V��O�9rk��5/PN�6�/y�N�'�*1՚�������r��Q��ɡ��e���|�֫`y���uʵ�@�T,���<�@Nt�9,��K�"{1Lrhv����h6K�.�0�Mrdq�)�p$�M2G���f�>e�Rk��/D6���Mʱ�ǟ��:�%���B���I�4�)��gQ�Ć�B'���ozKН?
P�(�_�6��Sg�L�g)=�e<�����9u�ΰSK������<������v�z2N��"�>�~���`+��5�7�ă��">J��a�#KȈ�SN�`�����1G�8���"�ƫ�Ġ�x��J���ѷ���D:�K�n7��T?먛͏r9_���b w�w5��Y��Z	�*�/�=�7._�F}��Q��]#��@��+B�d���T�������Q(�oC������K�/�柕n��Ҟ�׹����r�eS�?E�{��VH�JY�>�k��O��#��O!�ՙ�Q'���W�������tc	-�� }nz�2�9Z�����Y�Q�k��\��A���c�n8֡*������ק\��mv�r����R�X����y�_۶��Xt3��e�5i��>[B�8g���=��$���:&�s�y������>Rf�q>n׺���v4鹜�qry�=?w��n3����C���_A��?���? Q�ɪ�6a�;��j`�Ϲ���i���~3m�wb %��:�L�L���
�}��A��1�����K�C`9�O��o�@7�����=
o7��a� _P)��\���r xܿ Q"�$��>n��Sm�I��U_rf�8���{^�IJ�G繜��9�C�t-�$҅��b����W��A)5����(�!Q��?T�2��^<���#�D���=Sʻ9��m
U������K��f�S�dO̎^x>bKA&��X��O��b��`D�@G�M����{�FɌ�L? ���7,�a��6Cg�A���(Ec֍w',k�՟�,;��Wl����[tW+ �O���3љ�w���U��F���)]�]�8<��&��/���@e7�I�����Z�Zk{��v6�E���q��|�h�h����ģ��U2 �MI�:XE'�+����_�)
��aASi1�;�K+K�sy��g0�L��6ѫ�����3;h,�j>��D��<E�{�UD����q�4&�� ��l�}<���#�&q/��>ř���P
�ܩ�'Ğ�I�+6@�W[b|�FR������Z�>h��q�g�񼯇�ߝ�����b��Ɯ�^uݔ�/����g�Yb�%E^���:�R�-J��
X���Rn}��`���oC��9��ʧlE���d��K�O}��6Q�r\�9�7�+��P��포�B�ܯ���N�X��	����l�G���P(����l�J�����!�l9���H���*�\>{k�q��H��}AK��"��r+��?�Ky1������W���+XAbDc�f�#���/��J�[�bu��y�G1i�J)���
�yε7�wВL��2�����֤H���Z\Pbm�ë��-�5n��+��U)��-��6'�㐸T�Z�M�]Ƙ�_+��n|�a_��V%���6W�x!�n�*B��J��g,l��Ѡ)�k}�wCM�Cdq���Й�1�w�\|���$E��џ>9��/:8r#7P�ę�{v��f+'.���1H<��'���2g#֖�R���.��J�M�yf��>�DaASN�k�`80����L4����c���b��R�(-o�p_� ~ۙ�hL�+�g��S`������E߾�c���Im�vL(�`��{���81�N4��0"�lJp]�.!���l[��T:mE��M0`�5�\�&��mY�f��������ʡ�7�L�ۣH�:9#6��?�X"p����r������DG�cR��Vdis$��]�&*B��N�ɨ����h��K��ą�i��K��ˏ�5K��!d�e��;���=�p	Y׬UZ:�����Z �Ҧx�ꭅ8c��:#V� ��eA�y����W�k��A�;���F��'@ܦW�Jؗ�u��O&B�:��t00R?KA��6�j������!x�u���d�	�Έ�%c��d���Ʉa�~�4gjB>$J^+�x�'?H����%�C��A�ߕ��Lx���W=�_Ģ������!��\�G)"���s�T�s�����2,���PH�5$��)��4e�?����R�.W�q�j૗�~�]q�?�;B�|_��῜�}h���R�3b�̺A�|�e�+�4@�Z-��bD]b�I�������p��E�a�%�v���QM_�@�]�7���1�B����QN/�����D�.EZ��X�X^�!8\,x���|��S�<� h�G��Y+j�����|��������3�� �
�Ɗco�(f�����`K������"����l�M	�2���)��'�=�&��Jԓ#bC^*&oO �>�W��X��\��U�k?��Ά��Lř�������K]&�9R-С�&!��_���	��#�L��s��b�����lCM���%��Fd%�v,���nT+*��4{	���W#N0�>�'ę�PQzK��|gTS�ҿ�r<�*�(��4!��t� ]��@h���j����J(J=�H�R��{'t�#�����?�k�_�e��v���<�L��<��|M֡�XV�����<A��6��|�D�U���i��iH��[����-�3H����ne\��/E\�e$����?��_��}|U��v6l�VH`�5�ז1�Ӧ�ݒ�j��6�QB|�� � L.�,S#��Q�v`w!�ZI��5��U4=�&���c��J�~$k���Ti���@K���~��O�{e��sR�-��(���-�$Gzk������^�iO�;�)��DR\i]��`f���,EB��'��g�=�Uh�����V��SQ9����y�X��@,�iD: �$p�����*0E�����j�(��h0oq�2Ъ�9�����qcrw6��9�L7�&�9\���]�������(# 侽Z׫FI��9�����7?�z֏fx�֝ �0��y �����)v-np�?�yGJ�i̒�=���`���!1a7X�F�í��*���>v�'$Bs�� �����$F���-/z�THl+���ϭ�T�N�@��&�\b�-����_6G�D���=>���)�5u�_9�#>d���0A���(�/�^���j���y[�%pH��y�Y�GR� B�{�,?V��3�C��X׼�P�r c�q8ޝ������(kJ����i��VHI������hw�9�Mb�>��l�jN�Cg[�`���$��\�J�3[����D)�!�ͳ��u�����fq���1+q����8�EN$>��<�ڞ� �u��{L�_=�-G��G�F�J��iih ��7��w�
ĥ��6K���~��Y-���ě�3,1|�w��$��*qI��;�&[��j(��H�y�9S$i�S��� w7P�Ա2��&'�����}�ei�q���w�W��{Vlڃ��Hb�z��]<r�D��H����; z]�����v�>L�%:f�6�`�kޕd=1l3U�����F���9P��Ʌ��(>G�ˉ�_��+6�"*�d.S�{Z�c?��_!�,x�绶��=�hH�bJ�I��/b�����5brʯ_��R�_AN*��Ai9ֹ���x���V�ON�;������~
��l�_��=�{�׊�J/c̸�[���Q�@Y���v�(m�ܴ�RI&<|3u�2�;c?Ѝ�Ş<��~>lU����Á٣"^�Ie�9�
lC������P�#L���*�s���O�^�-}�D��H�D��S�fyhM��v#�͙��e[���h6�j�N@(�e?�?���3�;���wF1�40_\sV�joe���׉ ���}��9�{���Y�~��I^�2���/��|+�����j����ҙ��w^�1ryO���b�]Ӵb~{�|�yƺ��&�l͹����.�q����6�`<�A,����B7�$�4�1DV�H�S[�)��(}M����f_.sq���Щ�K�6���;*�]ju�'�������0&ѓ6�g��?��ҵ֍I��k���b���j��9H�0��?�}*
#�Easn&��E�'k�m��vJ�/��yu���R-L|��%JK��h�'�3L�j��:����'�P�ӧ)�p��i��ީ�%o}2�t�|>e���:h�8u�e�O��בݩ�W%~��_ݵ}gl�9�@���,V�wVP�ӌ��B���Qߟ�sA�	�3V
�}T؋L�}��H���V�5g��5i��Իb��\D�<!�ǌ�.����Q��n�k�>�_>�u+ɢ���&z�����׾4�Go�p�S��+`��j{v�FoEx�
J���a���1��ԊL���!hk���m��޼���g�e��Q����齻���%d��^�	zb��fb���_�G�s>p
�$����ck��ɬm��ú
WV��
�&G��"2O�T1~JOfW5M��ΊSc*@O��7����bؓl�12<Ŏ�0����!O%|�Q3���7ν]N~�4r�CԄ
�(���<�
��!ZI�7����E�s
�Д�ɮ/�5Cc����<DAN�:��U$���B^��	�����9ܚ�����[�1!]�A5˝�-�Ԫ���!���<)�j��2�K9�q][��ػ�+�K>s��ïK�C!G��.��db�@��#+A<֨�[������s8l�,7|��p�͛�:���񮢼��Rc;�Q g-VO���	g��ᚾl@�ȎSg�N���qP����`�-�U2(��Bxn���^�ZB���w=�I�t����8(��F�Galu�Y��\�҅ ��bP�E.��3���?.[Ⱦ��h�n��E(��6�{�U3��V���:F���U���L^���;�����>"�xD$�݈�Z�gD����n�l�p[:J����у�^���*E徕�//:s�;HK��&���ļ���yy������y�m�/��Χ�PC[Wb�猯u������H�#�g�T�y�E�Y�ce��<>W��:��5�Y�қ�"_	�����g����n����8�n�nK󕼛��*x��Ss۝ �~n!Bz�מ�6��-f[����[^�s�� eM��MǼ:��r=��@��F��s�~���j2廬�M�7��E�|&x]]'V^�����`v�>�B���I���V)�����2���I6f�l4=g��7*4a�� �>*~⺼�H�pIM6�-iFm3�����]0[��).pA�u_GAAM��P&©�T||�kH-4=�:NE��8�H
296����Z=~����^7-��u�~>����m�ys[�� ��|2���E��+O��kq㥵����b�N�V_�&�˷�r�˴S֬��ļ��ng�����WE=�\�rݼ���6�ƻX���=�|��#���K�Yd~S���{[fl��AȤi��;4��� ���Ҋ�.����Y��-�f!�e�z��������Dw��+�V�6!�>�|��xW�ڞ���B�aޜ�a=&fEҾ%�w��H�N\�
q)�s83��U���<ٵz&���:�*&C� ��I��T���wW��t8"$DY69|+M��w�辯���?7q���cZB� �ķ���F	���᧪������x�EQ]ѓMz��U)爛t�B�6N?A�ֽL�`C���w�_-��EP�3E��N�]M�H�q"D����HI{��3w�@m���jF�$�6�ZJ �B�yx��-�Vi]�O�<S�~�k��]�.�I�+���e�_v�����z��f�Q&��{(뉡p�+�s�X�����H��B����j�"5��|Zk��$�=����+=��?`4l�k��"����=3Qx4�ܘ;��Fn&]f�V���Q/D��z~գl�S]ct��ڠ~:�h�s�l�ב�Mzѵ��W<HSUiW���.��aH��O&�0U߸qRk�SM&�i-�yxńY6��˜O�5!�Y���<�(����E-��=�~��ˡ�j��a�5�����ƩU ����U�:C}vaf�Z����U�e����(�TWTjm�*���"
j]kڐ#B�Ć�V3k�^��U��wbv[�R���UҦ���b^!܄�xL)7=��<Q`!��9�9���g���&��ز���u����(l~�I��Oj:�*q�-C�x��[����d�ƅ/o�sh�
��m�C��^*���yB�b�ʑ��ؼ�`��B�\���?*��8�o�:�vU���gy�)����x"ڋ!Mc$���.��V����<�v2�mF	p�9�'�f����э,�vj
W�����5�6*�����ٻ^D�ϢۣD���&S�Pz�)vz�dy==�����2�a�5����M�:�������p���Xt6N�3G�0������c�>!�UI)z�X�~��YNs!���86�]����$UtK��3���*������6�\���+`�xU3�UQ��#=->FnU͒i�I��z�c&�҂�i=	�[�����i�ڿO�f]Ii=K1�[�D�A2b���S�]���"��
f��a�����Fs&��E�9�/�!��]&�����d�J�=����V�����>G������r1P�E�x�A��za�����(f���0*�F0^��c������l�sE�Rm�������Z�ΈL� 0�e���!�*�>�&�N�BG3#߉:���F�4�ÖP>a;�L~iɔ��u�lhk�UtWN]jdcFsT�̚e��`٧
�i��}�Hk'�'�v�)�0o��=���ꅽ� �; �5��9A%�-�3��C��!��OMY���)��՘�oÄ'M1d���j�>0�vǡ�FV����'JJ�7^�d�K��Y��Ĳ�d~Ď���t��w)����e{�l�=���w��,D�N]��V�A����Co&~2�����d�%��r%]�9�_A��RZd�yv�L�w�|Z�?��u��f�BP"(�Tm�6yS�s�,�t�!f�� �^���e.�5�ɰ�/B6MW�>#N�ڟϷ�Q��+�MNoǐ�<�p���;w)9�T��%�y�%�w�`j8c����Y�SȔI;�ku���ܪdh��'!�l�L{���F�:�<������4\��v��E,�;�݅�Cx�./�)��.�����iu�����i-6��j_�;n��g��_>re�oJX�K�27Z=�u����7m��ڊrǂ2[��:�p����id���@�D.)���o0��ZX��q� l�bTJxs5�FN�1D~;ʜ`��j_'!n��y����XH����2��qO�к;VD9��]{zr��z����T�:9����t��M�a�:����r&�I&����Q�����up�r�o̠;�x�茪r͢}���3t& �縶��Eܕ .RW�\j7#no�\a��v��E�v�yr,�˒.8��*_?ɬ��厏zsಭE�؛�ͳ���<\D�f"�<$~z��N���y��_��Ȅ��/'�
�X�ŝ��G���Ε�B7zu�����q���� ���AG=��`ŪƟN���Z}з&b�ѕ���[ZY�4� �i��Ui7��b��SB����\���O7��6�%JZܲ`�������ycD^X�90퓺%��3��@u{=4��*#3mְ>����Gh����)�Kq�f���ex��k@��r�5�2�~���"�eI���L�E	d�|#E�vee��&�����:aj�s��[q[����S^U���B�bEN�V4�v�a��\T]�3�L�߈/�jh4�H�Zv`�X�G����2�q�-��b���<����c�l��:.���L�h��N���K�x�!��2-�:P�)�$r�ʺ�)*q	�mu��XM@n0�2M��ݍK�)�\���f��y��{uP)�� +�{�d(�q�n�Y�BT�c�.�	��2<���lz�-P�}�Y�
,�P�p�j��q����	BH;�P�N_o+w��2��(�0`�d'�9�**���f�9�U�I0���@N9r��
�������7�l!6aT�9����Bp�ԟ�
@q�|�i�L�OL1Z����H��ۢ�r��3{���]��ʖƬ#��g&�DA�V+�"��{��1�	o�(_����T7����(��#���L�c����Π�O����:��hs�\+�jZS���u�����?9d/F��<�j��h���D��U�_kDܪ�v���L(E�o���5���֐�<����\�0��k_�ݔ~�o�df��|c*��&Ҵ/�t��'����+��9��:�'�eEy���.`���x;�F���0N�wI���1RW�c�W4,����	R����kgZ����D*ՙ��fɻ��c��GX:�^�͹���}BT:v���@Q��Z	��gdϣ�q�[�2����\��+�}���W�~�<j�*��N�$�@ԑo'y�!X�l�m��Ê�q�@2�5�"�����+\�E�9"�� _�#y�N�F&C��Gt}orѰ���D-�r���l��-���<����'=�P�eq���>�K\���(�S|A�7D����"$5h\�h�z>�N��?��S���ʂ��������^�$,K�Nȹ <��/Y�<˥�4r_tg��(&���I�0qd���"���i�
��g�{"�b�o���C.޷�~d��$��3����}`MG{ &�E�25����Ĉԭ��M l�����	Z�g��.ўrd�r�Ϩ�Ѻ�gg�ý#-�M����w<:�}��Q-�b\?���w�K���d��m�R��YJk(��e6��k����KxH܎^8{���3�[�i8��%×Ff꙲T"��x޺f��M���3@���$�����0h2]�G��+�#���a�v���I��Yқ���D�q��!S}'{x�ی��th�-*�ś�w����g��@�y��V��BL�e����.B ����V��"x��˜��] �+*'�a��M���*�����#���s�c�A���Ğ�~u���Y�ۼ�1��"��Q�ǂ*0�`�H6��%� ��𲎔�N�����?��ap���)��P�}��	����|-u�� ue�%��I1=j:8�~v���[�~d�T�*槣�c�EPO���X�L�n$�*4Z��o쳎o?
Q�T��|HA���ˍ�oϥ~�g�;��2q/�������\�_Ey�������P8�s�bɻ�ĝ�)�0&B(�E�z�ü+��-/?"#�E���[5a��%�}ZZ+ e"Doq�g���'Rm�U��*�����U�Gb$X	� �>�͔S;Y�`$��U祿��r <A�r2��u������#��̇9��W{���"�K`.Xfa[�U'ٜ��R��bh<��{���
R���*�* �L?>]��L:�Oy���Ot�^►1��b&(��*=G�6����2^~��s�VM������K�1�X�����|��0X��9�Ogz��@!ޜ�0IJ������M���u�}['h��ow&�_�hO�)��F�_�d��
r|k���O8ߪ����CF[�E�	�J���!��ʕ��Ǝ�/ɽ�������ukך�i���b,� ղ�pkB����?���x�tu�DЭW�PH��1'������S�R�$xxU(O|W�Ş��Db#i�����<���^,���Bo�"���HuA�2���#�i��F-YC�!���K}�.+A��P&¦�����)!'�ȡ>s�'9��ݥ�jNsO��QcC��5�eI�pO�◱�6���Q���`��	�rLaM���m�Ԁ��%��lw��Z��c)ϕ���y
L��h.7yz��Q*ɍ��S��Q��l�}�XIe��Y���ɩM ��i�e%�4�y�_���	r��LE��E��!j0���ɲ��)��S������`׆�Ǳ2ޥ������d�,��[��.�窘�J��7�߽���N#eRǢ��ɳ�8��>���	z�q0@}����j]��l�t>�)!_(VX	ݺv��V�4E[�N������3 �������$_�.��"j�����Jd6^��&�~�I���I8�H@$GT�&�bˆ�Id̲(6]����3m�[�,(,I4a������DT�k�?�\J���=��(�K%�:Y�H3�u2r}��h�׼
Q��u��m� �82"����%��L���%M�����Ċ8T��Ha}���[U�dX�>.�6+��'��tN�ʖO�ٰ�4��ƹ�NJsEa��/��~&��W�������L���zD�!�-i��1?�c7o�aR���:�SGg���pY��C+߰N��4���m����CZ'��N�I܏�_��4�i�C�"�a��Ä�$��Оqn���Yg�m��Z�̺�����'�{�V�+��f���{.M�7ʷ�G���135}^+��B�z��o��ڠ�Bo2g{�>jwb$��Q'�̐��p �7j��PX���[p��r�Aw�5e��M��W'���������b�1�n)^[F7��x ��:�����/iڰ������k�o����A-�\��Ǳ��؋�;�ͷ�pK��z/{wk�N!���V��Ҹ��u)i�x!m�������A_�F!s����?�?���_����G�/9S���ҭ'���8�������N���H1���?\��7�s?�$��_a�}T�����\b�l�255��7f��
`y^�N~��g#�m��r��|�;]mdĠ��myy�����NNN+�!��1��k+�h�����Pt��eT5���P�/���b���/��?�1m���������_�/���b���/���O���˿p��RCE[9�����PK   F�X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   F�X'�Sz�  m  /   images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.png�WWP�E �$�.��(U��TAz/�J�.AzI(FRT:"A@� ����P�j�b@�����>���93;g��즚�2�x@  �Y_O�좺_���"�\� ^`��m p����ma~r�ޱ	5�E�{ P(����o��K��L@���-u �対�-��|r0�����|{22SԈm�����J0��d�]��r�2�~�:>������OT��9tW���,&Z��IB)����Me�iQﭹ/��G�����vѩ�6J	{NԜ��O��:(s$|�T��a�k�W�jjn�cX��e�!|�1��/><=�Q�����uu	Z��y˜��{����Z�xc��8ЮP!�Pݏ����]��J�x�nUz��tY�KD[N/�!�n!h�t�-�)�ZT����HXQھb���3f����cn��r��:����?L����m�?����#"�_B>������+ń�N�O�	'�a�!S̡�ɳ.?�K�+糮_�1zU.D��R��s��LM>������IZ�Uy��N�ʻZ�=^1����&��/�j�{~�B�6�$.��h�	b���K�
�Nv�5<�5U:�ش��ґ��]|dӏ`U�]g9N+`��&\g#�&0Ii�~Wi��qF��G��Z�ɻ�<��=F#P��{�q �?�(/M�fś��&����ؖ@��9�C�L�r�KV�%���gV3)"�r���9���A�1��K����&�̑~G�ZS��`����z�@������2\c�)��u���fY�U���J��������t����N§��r��n�DT�ם��I�4ca{�4�R�/g^�Z΀����*�]����6��H����4�����ђchw�n��In�9�6s�kž���s�_�q*�8lJl�$�B��J�^!���g��YGTW��{�Y�Kv@�~C��N��p������:F�I$�y/���=��}e���!7	a�y_�,D!����\~��G���1K���۽��P�1�^���K��]/��gi:)/DT��ձ�W��4�e�����׻�TP���N�Ĵ�{�|�~+� ȿ��TfT��_v�]z6\4�^�(�/�?+r�^�-�R\+�d�߮��`vͫ��I����R�2���#�:���\���/����2~�ޞ�6�OT��A+��U4 �{��V�n�L�9]	&u�Ê�ʁq�c�IW7F���&�ڿ����:�}؆��٣��C�ܚԟ[k�&��>4/irƛ#r;���?��!�:�Q�n��j��p<�@B�0�?��`tty�j��~�✫~����]�͡����}�`洴z�hw�S@'2f  ��!=�7��r�\�pW�쨏����C�����xI�����TIΨ���Q
B��������������D٘!��|�^���t/v��_��M�����-9
�ںmE�m�K�
��{�(��yw��2'�y�4)K�	�WN�4{~G�"��p�^T��W��z\O�g�Җ��N��?��g�g�a6j������o{��xq�VD���r<Q�R�.Fw�����X5�͑�wQ�d�@�ݕ�0(�!`�5�6�8�.HלI96�<��X*����AoV��W_������ɼ|����.$��ڎi���J��Σ��j?��1��Ս��tƛ�|�;N1b��3c	e�~ͭ�W3ɾ9�2	4�';+�~1?מ�\np�E���@�9���4��V	b[>tҗ�Ψ�\n�O�G���B�$�ܯ��l����bH���r�(kDJ��o��������50qu%�Q&�l��q
ah��B$@��T�>3�=�KR�a|D,�'�RD�7[w��p�e�	m�`#6�-�z��/�R��I�A�S�ݥ6������H�G������׸�<Ի�}͒A��)��?iS'۹�dq�@0�p���s�uD�EJ�~=��[����\���Ű�˺U�Q�>�N=�)ߡ��h����Q�C�t�V�g4���5".TkN�l[���?`�z �"�����9�� ;41�r�0Zv��͝�9��E����hth��kK��iea�a'v�/IT����"�R�aQ�2��Z7�M�(�@�8qf<	҉x;W�+�\l����?��߫�å��^-MW��<������:�[��(�Q���h��6@�2zP]A<,��3���F��[��~��6͂�J>
өQ�Лw��z����	8��/���M�W�n�=�ѩ鮎(�O��N���'�bSK���%��C�L��M*sޞ�嚖?Js6�.Hz#�o`�]�k��Ӑ�J�}�gA������N��[��j�
���&�u�Z���,4K�:&��V����W�����w����'dӧT(��ϏvpI�1"���ԥ�[�N�C����l^!����d��[N�\�������y7�s�������!/�B�'S筱d��(
�f�Lc�� �ϕVG�֜�y����Y�W=X���C=O�x�?�}�Ͼ�T8Ab���'�r�}����+n����o�8�n���Q�8M�ubC��S-Wׇ��Y�Y�^h��K�[���y'�>0B

�U�d��� �.Eo���v�[W���
��mYe��>=Gc�ְ�36ꍽ�J=�U1eR�ѲoR5�q�DL���>.o�ps���t��&�V$�P���s��H�3s����t���kJw�Ɠ �K��YK'}4�����N�; n������`��~�Py��S>�_}�ff���{-��h�YwaPg���UAt����#�c@A�τA�5G`��{� �'an�')�,�8��&���2�>*BaW�c�C�t�5�0m�niz���M�c��I�0+�Ԭ֢7��q��H��d;�s�~��q� ������83�{�h/�#��nC��H�߳���v��M.�����l�ýM����,{�	�!b:@��LN`�gIZ�I���]�MK��͚o�/ܨu?�Sj��Wbo�	���ԠJ�1/f�S|����ۆ����VL�
��d'�ߩ�y��
��:n�P&)����fb ����T��>�W�Ŋp�/��>��R긥��O�9���W�J�W;�Nff��^8%�Ƿ��R%Ґ��&�YBi��3����a�����r{t?�)��⺜�D>��avN9��/:G�
]���i�alMzy唣���>2=v��"�DD����MG8�IYfڑ@:��?X�:��[t�<�MT��h�v#�lk�.��k��j�i79N�n-N�Չ@�ۇ��%
���!ˇ��&�M�i`,���/���;q�t�쩉�%��v���^���`5��o�½���gnΓ���W��������5������+ŗ#S�k�#�g,=(�.o��?~�8�~PdbM��z�S�Q���i�v�o�ք#���Y|�n���xSS)P��Kq�1��J0D����[Z��u`��Gmo�$}�:����8	y�;���7{�?Lg�w[��w������__��;�1A���M|��gJ$[ܣ��w��{��M��&�-VL�FB@�L������5��_/D��{9�|e��\�s�i|mx�S��9i��X�z���R��%�sہ� �1�l�]��5�^� ����ɲ�5Y9�9�M�G�V�׹�{����Yc���7i#���T�S���Ų?�D��^�ˌ{>~�!��82T�;����ਊecС��D�S���W��X��L�/PK   F�Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   F�X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   F�X�-��_
  �U     jsons/user_defined.json�[o�8ǿ��}�Ś.�I�ɠM�$�`Q(�J�:�G��v���KIΕ"Mo�3؅�P8��;y��^�o����L��땩�L^�&�Φ�M�*�Ҿ�p���:i?�������'����~������7�z����n�uU���/ҺJ��������������^�+3���TQ�s�9���F ͵��RR����UZ˦o����"�K��08��D$4@��(�3(E2_���{�oIK�������ލ��β(�˼��}����b�\���vĔ�9�y�~^ݶ�1��wֺ,~[�&���ES֞���ժh[��X�+�08C�}�X��Ǫ�_��5����B'������ћ��a*r�t����8,v�,
{~tqt��ˣ��x�ԅ�((��2�˔Q̷'�^(w�껡b�:>�B��Q�}�e*�����L��~WT8�����j
�9���I��(����u���\�����p���s?����}ᇺ�"(*�PWP$����
��:�_Qȕ��~��v5E"��E�]Q�H�G~UaWU$R �/+�ʊD* �u�]]u=��V�!F�.��Ѯ��!�B�W��~��h$�W�m@i$-_]��zñh19���my����b��_�d@�0�l���!�MŢ�mu =��D$N���92��b��&�!�@��N;�~�@�	�]E�X��0y���U�
�X��0y���Պ����M�8��&m"����y�$#F��X,��38�ːL�H,:�C:0��q��|��"D(���SW��qC�u��"����d�6M���Z6P��T��ٚԠ-�EP���Ԡ-�Gy��Ԡ-UDP��;6P~�TA�W�l��l�*����s3ݎ�@��a��I`�
��#���y���:$��}����q��P�ȸGa(Bb�?d�#1�12��P��p`�<"C*Á!�,"-e�+2
�;+pWc5&+�gCXG��
�y�p�Qc��uJ��1Y��:'\}uԘ��_E��:jLV���.
c�B`�\u�ؘ�/W]=6&+�#���1�����ȤG`QY�?dң����2�XTV���h,*+��LzD�C�QYdV��m�^��׷Em2ki������b�M���^�6gӲ߯�Y����z��v��A��(��f�o#�nO˃�fyo�ݱ�*VE�0��j�ۺ3��Ҷw골�u��f]����~��L��(Ҫ���SD��* B9�:C@g�Lf�d8�D�;wj�T�)���dI7�ڼ�R��W_ؗ�_S�~4�p>���� \�C:�i��zU�E:�0�jo��)��r�n�{�H�m�QL��H�Q�b��"�c��{�*Qki �	� ����X���f���?s�h��]~5Ǌ�KN�m�L�����#��-��W;l�˖n�z���ty~�v���i=���t�	�~8�� �n ����t�������J�?=$\,u��ͺ|� 7J)(f�Y�<��(	KlV�R�1a�	cLc�Ƙ0Ƅ1&�	1�J����F�7USՓۢ�8�rM����,6tw�ۻ�JRb�K�d2(5
d9�@Ƙ@8Q�(Xj�*��v*�&�ٴg�s*QDxPs;���Nt���}��[�k����$,~8=���I�Ռ[>�x�E_���
;?}!�?),����\ "�'W6�XoF��
3*lTب�Qa��F��
6*lT�Uaﰒ'�ÃI/��.>���2��f��L���	�m{U(�3H�J{��њ�2I���V����$�vJ
i�i-s��x赜@"�Aθ��f(�8���\���$f5��V�*��]���#�f��9�
mY�9��r'!��)�6X����-?�T��'��1T�l0Rw�=C|���w��F�1Lq,>xnv`-M��*����<(|NTlF�#A�sj[z߿9>p����p%Bۖ���Y/�Ԉ�/�g+�@�u%��9�G'����g�x��Gyo��!�=iȿB8p��f$$1e3�a;(r��ZK?��)��$w4�����$�S=��N��z�?�=��)�}W1m��$�O��hc��`!�IO	�ނ�;X<�;��@?�J�`!�����)~�_�d1ux~l�̿��:|s^%U�2��KE�� i���k�4�BOk���v��,�4�UD,�@�L��N5��/Qvz�s#S�P�UeK��C�C��AyFAµ�e�<�$չI������i�����w�ml� ������1'>�n��Mφв�\���-�FI�I�M1�#3�)2v�k�9R ���$G���Ѡ獾5���[�o������7�#���^ٶWۘĜ&h��PB5� �r�)�<֟��:M3�����F L��<Mr�g��t�����.��}o>t�M�Y��Et���!weLc�4���2�{V�-��"�4i��Ɋ�O�o�t߾{C��l,�-VJO�i�(�w�l����xv�ݗ5��t��O�u�.3+��q���7ݿ�{�.u��Ў����VA�	;��l.��ͣ��� �!պ.L=91���<�3N8����֧i���F ��l�d���G�^���<�y���Qϣ�G=��z��ǿPK   F�X��=Qb  �L            ��    cirkitFile.jsonPK   F�X����7  �  /           ���  images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   F�Xs!��}  {�  /           ��0  images/330d02b8-4530-4fd4-b6ae-26fc03cafecf.pngPK   F�X����(w  +�  /           ��G�  images/42266fcd-641e-4cfa-a619-b442e1b7bf10.pngPK   F�X+���  D�  /           ���% images/5cebb09a-e86f-4cb2-800e-22da09d26481.pngPK   F�X�IM��  � /           ���� images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK   F�X����H   C   /           ��J� images/8e6e9996-4250-48fd-a42c-980e5b13088a.pngPK   F�X�&�}[  y`  /           ���� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   F�X��) oj /           ���% images/9b962a8e-14b5-4317-8666-1954827ef6fe.pngPK   F�X`$} [ /           ��O
 images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK   F�X'�Sz�  m  /           ��y� images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.pngPK   F�Xp>r�  �  /           ���� images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK   F�X�+�s;  z;  /           ���� images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK   F�X�-��_
  �U             ���5 jsons/user_defined.jsonPK      �  T@   