PK   O��X���  պ     cirkitFile.json�]Ko#7�+�U-��$}�f�!;��lC�;��F��d�ߗlI-��R�E�9�&�X,V��Ţ���>�ռX�v��֛�z5��r:������S2�<-V��z�k�=}��}�'�?�lR�?=�Wv���<E�W	W�MD�T�e�$y�)�ª2���������)�;�u��Xg!*Y�2O(�<*5I���s�����S6A-PCs��7i)���u׸�	W,ܑx�H�S��/���أH�Q$�(~�?����[$��?��KQj[`�6S��%jl�e��	m]i)M2mK����R��T�p�Ҝ��/Ƈ�M#W)-+���**����X&Z�D��h[d��)fd��F6$5�$���u�J�(D�K^έL�9��<'�,�y�֙P��E��b�ZU���gF�!vX#����SKY��eB�\'��g0N�$K��jJ����tH��FF�t����m0�{H��6&n[�4
�w�;�S���:�T�Af�Vi��C!����R+PO36�G
�4�B�M)���6ᔸ�3�0�,��BK.���2MC6��R�=Dj��:�1�6F�D+�\+�,�6�L�i���y��B���8"7���e���.U�/���#��`��!�l��
�F�I(�Csm+��UN`��(+���DU&�Z���mpd`gD��h��3���3;#f;������P�OTl�9���������X/�5�e�w�� �]��{.i�YZ ���,�U�EFy�4
������A]$��A/�_��q��A0�a�4�i�8(f�tp�8(fqP�⠘5(.�.L�a�G���B�8(f�Jr�Q!��bI�^B�(�#��?��A�r��T~.{�R)*5�T��O\.�`h�=��.�&�~�*s�aC�H�.9��,�y�q>������:�>�RД���M���NД�y�M_�W��T��y����4Ex~^�)���M��WVД�S�m��,��T.;CK	I�8h�(z�\C�9����i��c�e�Ͷ�eY��m�-�Y<���ED�"�pI�pQQ��(\L�Eo��8�q�K� ��A0�a�4�i�8(f�tp�8(fqP�⠘�A1��b��"��Y<��gY�\."�e�s��_p���"z�Y<�8ؽ�G��,�ā�e?�e��&�/��,����gY�\.�β�\��e�s��F�,��EY�Y<�����,x.���e�s9�������vW�2_��ON�,j��?-���j��K[O��1R��|�b��0@�\t��yf̩�TF�9�����@#�1$���4�7xfp�z�g�G�6��8:��EטkB�`3�s�Q�N`l`��`���Р�&PQj��!�.t�:{RJZ�<M43¹�&F��r�X��+sfc�z3T�3r@�����@�kXi��b���[<5���#y<�����"�lU��N�7���!^#P8+�k��@�gx��/ 2�8+�k�x�!��f Y�l���v4θ�.��gx��/:�8+«� x	��^tDAl`�#2>9+�k�)x��s#�ˇ�:F�{� ��GK���^ �>��7ۉ��1�Ї��*�J {�8���6���Ū�.n�^W�����yQb��ȒcL����+H�b.��!;�$��Rd�쯑�]hxb�I� m
�P��C��!��b�ȰHdhM�E"�"�a�ȰHlJ{�9���k�{���S�A�3C�0/��
���0�cِƥ��� ��.	ۇ;�`g44���t���:�td�.�|C���Vx�q�&GKGa�^�C�-����Rd���$�6'�8��.�g�U�=v�����-��\��;p%3l��%�=v�m�m��Ge7"]@�˞#��.����а�WD�VB���#�E��A���� ���A?c~M��z�<����[��bo�bm�ScR;�(�����9�������`�kx���`��=�S��܂�M�����
�Ƅ��㘮D�v:@�^�@uE�N�v�t��� P�tpH~�xe�������7�Pq��CU��X\��PU�^���0Tto�VL��J�f!�U��o�~�"��˸_��|�G������"�k�W�c|}�͆a�z?��A�ޔ��0L��`��0L'�^j��10LF��s��D0�e�^}��W0P�/��}������r��.]o�� �_v�7�Rz-t�D�Ml�ĆM|�ćMb�$�Mr�$�M�)6�}�6�}�6�}�4��l��t�v:��A�A�BB�3B3��"��r��6+�uV���j=_.6۝niѱ�>����k�чz�d����P�K�z��6/��R̸!�8�SN��i�2!��ѩ�����EUT����asq�͒�	�1�u�7qg+�/�[��o�U�c����u�p\����z��ǭg�����?�=�j&;H��T>N�b3~�B��tF�:p�fd���L�!�Dh���dK��C�Yzʊ��'���S>�b�s1Bߓғ���g�1�Vbt��e [�2x������9�����/7�┐���� ����I�"�q��ƥez�Ӷ�!U��z�e��n;�|A���-�?o��ź�g'�;-2��'��V�~7;�Ͷ^�~u�i�}�����s�|�}��;�˹=�N�L�o���/�W�p|'wU��X׸��/��"_������yQ[�ͷ��u�S�z��b�\��� �d'����:_o#H�U~��U#S�ε[z-�G�*;j�tP�t�TY���8s�V��M[�]�^�����joi���Kqh�
bf��0�(�����T��O �|���Iy�\��Ҍ0�G\"t�C���=!:��(���	eC��̤B3=��S��Ӽz/���qr�5=��4@H5�Owؑ^65Sʤ�!d�AѲ)g�*rx��3g�����Ma�Ҽ3qG�+1��oR�՞P놐O��-�vS%:7B(�*=<n�N�DT����ia!B�0�R���<��5�O�K(�
���SV����*�rbn�pA%�ӄ:%X��G�S�$x��������$e�ʤ�RQ���30�ʽ�u���@3QoƦ=���}E��Q#�ӲSFf$u~;`����(ȑJ�sP}S�|�J83�&��� ������A:���4]�п�)B���Ot��zӛ@t
��H@�Ƈ���Ѩ��JQ}�R257U2�cX�u�b��H1�ʃ�y8�Ci�|^�7%�T+,�T8����'H�i��_���n���'7,Ѭ���)R�cg���~�t�������p3ĥ�/���	J�k��0?"���F��ݿ��죋v��MfTR VȻ�I�=�Q����TҸ���a�v�h��'���J�r
�V���ÙWF.h�c�}���C�������yU6�j�v�}�,z�ּ��$�ϸr�7���,��G�B9�����?�&��>uQ�̅��۱��}���+���-�ks�j������~���F��a�|{������>�����Y���~X�ޕMӋ+KfvU�e+4iX�ٗ�c����3�tO��j�!�~lx}}xx��#�����s�!l��w���f���Ҽُ�'�6TB4�"7������$�(�㷇�7��.0v/�V��+D��`����ej��|���Q��X�sP���C@`���@��o��q�h `\!ݕ��t���<]ͤs�
���9\�2�ȉ�2`�V�Ye�m��]��]�pјPA_B�#K�io �񬢋�>�d���|�]#ۛB�9!=�gsT:\�M���@D������`ճo�����O���@m��^"����Pp�ʗA��U3_�h p\!ݕ�89j���=mhWs�jd�;z	Hu�z�P�ΈC���U��	|��M�+�8����I�,��޼SgD\�k
\�X��"�"��]�|	�@gDXrX��,����������G2/[��{����H[tн��_!d���]�8��c6��5�EXJ��$�R^7���o
]�+���Nw�	�m-����.���_�E(�R���h�A��"�^���Kw���z�g��X
����]ǋ�wc�^u���������푍�[�A8��%)�*k
3������-��B����Sm<?Mw3p�K�Q)-z��u�����*s�hqO��]��Z����%�hH6��i�YZ�L��+��+z�l���dA�w���+g�z���J:�{Q{բoQzZh@R	�U�$��vD��> q����� ~�T���)����38���g@6�����TQa�!��}�Fp|x�|/�@�dEǏ�Td���]t����Y�C��d!�+Ն1C26�T\�S���1u������C��w��*��\��0���H@]#[�S�e�������Q��z�K�T���:+�%��[�|��/A^,������r3����4,�g���s��n����~���y��|������{�)��Ӿhz���PK   O��X ���s� �� /   images/25c207d7-bd9a-49b1-b471-35e2df67a92a.png��csfMۅ�ؚL�m��Ęضm'WlOl۶��m�zs?������zwUW��{�u�3\^N   HJ�(  �  h64����|Y�� c'��  ���$Q#�  __�"��n��0��j�d�9��ʁ�F��V�#u7�5�ƣn��50��n�?�cm$�?���.��=~����t��&a�̀����3x��e#d���I��H��+j��ʼ�W���\������U�|Y����1J���0j<K��=���&�9�7����<��K�QA��-B!�[d��p�+e�c�n����뀿��T��!?d�� *8�[����_q?��LPW��'���Yx�w`W��X��ꈴw~��E��m6�Q��V�ņ�Wߌ�m����x(≥��\�Q3����ʻ�ӌ��f�p	v�AU�rn���ŷ�%�1�)���'��%a�sO��U���rӶӹ�p��"��w�ʽױ�{xj�㋼4�(��4���n��c�7eu�P�K��p���hv��{�Z�����q'���20}�_gk�3�F'9_����.*[G�6��j)IH9�X|nR�:�?��0!�@��G���B��i��M�R '	3���Elh�X]	�qӢ�����+����&jqy(>��=���������Ų�1"�����1�~��%�]0���N5>,�Oǩ�K�\���`n �2���P����b��m��[8��X�3��f&8����4]���UH<��xa+������0Ӈ�5e�e�B��Is��>�����AT���W�mK\��}=C��ie�)�>��ee+aM|�i�K=`���OrƵ���O>*$:9ݭ8����)!l��g�S`�:U��j�,�균����o/<KNj܊�}����t��� x[�nɤ�Zr�[a�}{�b�q'(��W���O0z�n�0��� ����tᗵ�B��
4ɑx\�^9"��:}�_��IH:)��۽B�{o:sN��u��XZ:o<��4����׾��I�0�M0���B|�k�y���0��p�<����X?|�g��T����&��9k��}�lb�F����d�t��2�;T��v��C���`U�:�8w[-#O%>��N![��}5O)�e۪�-'f��4*=���ƺ�~O<���X�����(�1T 4p͏���2v�*�icd�x�S�����U���|��k��z���K,�Z�4����q���_�Jqk�������6=��c��{�
=\D�fƃ��p;�u���e<D�$���7��\E� U�6�ll��-l{Y���DG���ц���@�Q�%�o��z�hNOd OlVw\��W*��B��NF�A�~��qv��h�����ĺ�px��L}n^r�>��RC.�֏���l>|�!lZsI?J�rn2||s�jlo:?j|� ��g��2%_��v�|li$(�7�J�\�6���6��z��~�|��n�9��W{_X�J��9����;k����,�Y꼚i�;�؈����s�&5�O��=��L)2dx��ϑv�Kk��+�>!��d��W��?r+����
��L`gQa:a�� SYֵ����b&m�D�0L���V'\D� 7�T|T
����J/����%�'v�xڅQ�G�I��d�"]����}4��}�c�}��X�Ք��(��]�E^�D]��f�V�|a�충g�#��^��F��m�mg��1����Y�G�����}���ږ������˴�'�c7��c�9Ρ��H�����^ T�q�����
�h}�݄ł�j�ȅ�TiT`M�U��&Z��r�;e�1�*��{�^@j�#% �ψ'�$wcT�l�)9,߻��L�'�"i�K�D �Om��ǝ�j�l���r��`��[ru˰|���g����\�Q�y��cQ*
�3�_��V}u�Y������-"��4���������J�h4bb�r������f�-S��e��&�46hW<��u_g�����M!�E5�c)�T�t����NOx.��1�YL��������܂�� ��V(0�6F�
�K�n�Ov/�X�cPCP�rrb�u���[��l����1H;nE?#a��s��*��������q��ULQ-s'������y����rСsr>�B#�uUK��i�}~ֈ�?N�B��πgN�u?dd-"�%���̥��[A6%W	C�	�����Cm�	�/��Ⓨ�Z���5v��#��9�v�7_��&0�i�2b�bNP1��M<`�v%��>�!4~��9|�'�n�p?���T�$k�~�/�Q�L��v���G�� �VK�����e��*�c�S&ډf�Q�F���.��iZ	[������+#���Fn7���|����.��w�^7��ziM@-G�W=�'���D�?�& ,�uMu	�q�v��>}L�|���6\�>z�|��=�Z��݊�����n�?w������m���3�Uv��)3\	���t�՞��Ѥ���d��N$!#��TvO�9�JP����F��E�G��w��V >�!7����y&п똌Ҝ� 1u�v���EDm]qL2Z����揾���3|V�U�m�Ax�ɡZ�<�%�<�R��d۾�b�p���W����*[�4u�S@����Ll;!"H;/��.d���b m���ֽ-*؋��W|9<�cL���A����H�p�v��Qkc��[�t�����4a�n�_.�6k4Ń�6NZ�����w�Ӏ�j�I*��]YD�G ܓȗ�	LO3Z13i�oJA��-�����MX~?7b�aW�u��i:���.��<ls���U����y4���'���B�vy�n��������7�P�bP�3W�}�[�K�-
3G��z�Q���V=��|56-Ż5:�I%D����1�I��Oc;���4����!Մ��a��XBWW��(ˠ�I|�siq��gkcc\KK�R5avV�T����i1B�T�PЎ�Bs���z��ζ����Tp� ��J�|�PK��J�gX1��h'V͞A+	t�u���W�k�ழ~����I�,��%K5��ړ�F�+���U�+���\{٧Y��p�O�����	�F{5⎊sv�gG���э�&�~7���|5zle�k�g$M(�{J��YRu�	F0�d��`5�*n-�.��:]�dY�K�X�`�U�?�B�E�����<��yV�h�U���X���XM�e��dI��rz�����O<$�rjk!���Wi0�1@cu�]*+t�u�x�d8?���؁�Mõ�z�U��w��{1�t�]�؀vC�o���kʒޖY��ԓKOSk��[떸�ʴ�M��$�PH�B��SI��/�<?�޲��w�ƀ����6[�_U�]qk8	���P�wq��k�[��½�Sv7z�Ǟҍ��q��Qp��$���g�d����Y��3u��鱦�4�T��gDY�����nL��cy�Ƥi�C�U��]���2r���1TeeM���G�pz�^i�%o����3ꅣ
��@"�|L�W���E�Q'�f�N����81qpp�}�=u�Y�>�����gq��w]u�d�v�z~}~xs�O�0vi�S��vd�/��xv>mjv��|O[7�̪�!��wE1f�Ē����ڱ<�����*
��+�A�sA�յ����R��Q8��d3!���s?�21"FE,���1����H��FbV�+T�~5��(�^Ey���ў�33B�Js��Єܿ5lR����gw�;N�A�$M0<x���
��4-��Q����Kͦ�ߝ+U���&�m���&R� 3�Ӕ�2�-�.�����W��f���$�"Y������"��݁� =�;��I>�}(F ~�!+$$�c���ʴ�j���u��q��j�p(,//�,oM����oʖ����ߌK��lq�!��"U8��E�C�n�~�B�i,5�z�C��X��m�^��럣`LP���_�%�/��9|ԡ:�v�U�?8qp��BkW���\��e�����>n[Z��5'��S����Ҥ[����.���rqݴ��S��m�?�N�Z-V��:��5`ٓ/�,oA��4���wƨVW:U4����cFk�"ۏ�C1n��y��e�h��Y����t���hs��OEL�����ZRjA)��cӰ�����~�uf$}�[8�T�m��P��>9?g���I {؅F��dm�a�c�4�N[���+�%�|dB��L� �͑u�9f�֝�����Vtr��ӓϣ��4ԁ���o����i)�U��3��*�Z�z�3����U�dǴ	9>4d9֑?�o�L%�ڎ(Z���ɺ����W,�\��Έ�_L��g��/��4�&_�7��ӌ�܀�β�@�a7#+������5�9���7\]]�{���:��|�u���|?_�����^��d֢m�kvޖ�]7���{�|j��<Jx���Q�q�^&���XV�RљH'�)IOCԣm�GdQwE����4�Х`���l�5���s?��2�q��$��w~���5��Xż)~��m�!u8��/$�TFu�qx�o �3�U*D1�jPf�#��Q�"K�<u�߀�q�� �>̮�;�c�u���B�.�4-S�萍
'���ς�c�qvj�vm�aw=��Udnԓ�̈́3)c�D��ڛ�xa�Yq�ŷ��,��n�>u��2ʸ5;IL4�L4�j�9�(-�x^X�l�w�LFDMO���e��&d�6���,�����}J�G�>t�:0jy<���iW��^��pMN�}D�5��S��6r��s�;:�����3i���k#CˉM=��2j�����	��Efv�j�<鸍�O����wX�V/�z��X� �� ʹ��Ҟ�S;�l�.CG^~�m!J�O�V�^��!z���&���H �u�Oz��Z��o�����0�^$�#)�:A�;$����Y��0���8�r��<)���iM�r�S���Ӥ��2}��.x��������
��K�e?���'��Ξ}83^��xz�mga�vj?�F �i�m���o\li+�}�a��^?q�c�uы��>��c| زj��=a<c��T�[���e#1�O���V�X�75gP��b���� �8=;�T	C����f`��;E�S��.�����r.�2N_�6�_�C�_�
�`!}������xR��H�ӂL��gT�b��>.�h���{b�Z��&R1�t�|lso� �?��>��C7*Z�O�p�	.G����a���#L�F��Go˚�:�Y(s�kxXvx]���]����ܦ�!Y~|���{�Xk�YF<�V-�J�*ǉ%&6�i��������mN�'ot�?��5�т��Ƈ��,�^�^�����ٔcImQ�Ah���Qm��0'������Lo!����E����/E}��v�z52%��RS~���g���"G/�j<*<�L#.��䤓���䝴{mja��o�O�n�l5�,ЛB˰�@\i0O��I������h�c x��)��$��\����?���I�vqro�C8�Ä�c�Nf�\��TS�|e�UC��.7�|+|�5
���3E�5�H�I%�"9�N2�j6�zX�lZ}�<�j2m�S�F�����6��'����uT���I�ک�ge��(��1lC��M#C��JN���e�f�_�OJ&���{�韔�Ih���Vc�y��i�ꔀ����I��J=���n�]���ݮ��g�6�Qna}��k��<&����s�د�h�@�Ql���ʼj�9ʍ;I����z;�K�r��F'���;V��,�#�����2��ˎ� �CiA�6D)؟f��FZ���	��'�V����q��\\a�E�9�&T8�_j&�B�����6�^����Q%s�-����e�F�ލH�G���O}�9U3��c���-��չ��`2�<d^�F �L�j���*U>��Y9��� ;�l�8~p�-�^o����F>~3���|8%ι��WW��ҫX�t���%� M��!���J�AZ�(�����0�_sCݩ#��T.QȦ f?�OcUA���Hw+�ι�W����*M��Ad�K���jH~+�aQ�G9f���!��N����D�`���e�Y��|��%�Q�d��
n�>\Y
�J�AY|���]�п�U�_��G����m���kX,���!�{�����&_��@�$�Μ0l�њ��eSS�c�GN���.��!e�~���c�����:��{Q�"��G���V����w�M[���uk:������!�NV>O!k��O�4B)�?���߲?����%�@Jg�����fU�62��(QT�\;�r%���MЉ�P�28[(���-P��S�;����Ȩ��L}i�Y^S�	Ɔ�J$[I�V����+1`�^|� ���L�Lؤ󹬓ެ�	W�?c��g�Oy��Zm¶Nߪ;��wB�BР�����/�Q?΃�J14�5h�~sA���X�
��e��Ƭ{�VT���9����\ƫ#�v�r����_�h�a�7���i�J�ƎE���FU�-�L)�9�
k/�Ǫ�.>�U{�y�� �ޞ� �o>$�����d����P��5K�1g��2ef ��NjE=�
.�5�MIi��ۃ������)��{�CM$;d�}r�@�w���xi�ʂY3�A����@*�#E�"W�&�b5�y��D�f|R�>m��I*{�b\<�]U�*%�VR��bV�g��_x�]k�"�@���@5�� U�q6!+�%	ۧ/,=�D�|�%���z\!_'^4Q�j�>�c%\(����.=�ǡ10�n[ˁss�Oo+�X��f�$hƤ�������U��5��|��M�V7ý�	�p#R?�ߕ���t'!i���p
���u�?G��S���j��S�B�q�zd@�����f[��a�HQb���_C3��'2�����+X���ze�����'$XiK���ďf�a��z-��}&]��ύ��P���~Wb��̓�hT�q�J7#�?'ޒ�'U�x�4lپ�$ʁZ0���<{1Z�z�s~p/o�z���NL!��6��q�\����E�����2 �n|3\d��d��O&��]|�A��Iqο�b��^�u<���"��?f+�h�c0�=Z��]B������9��ٱɎͶ�h�\k�*��?��Kg]~<��w��-�p��~�郘�C���.mêyq'��� �矒~-��<7��#q0���I���*]�a2�����$����T�M��Ha�H}��Ր�WjvL���p15�Ux
���&M~G�칇��Q�(]Q��I(�˴�_y}�[.7�]�D��|�,'�� ��+�}? ���S��=��n��|�L������s4��)�**�����7����ͤvv�����8��f�.��gF�%Nh�,<뤠�%H�J�rH�$d�
�V}��M�+gn����ϣe�ӇW�C�� ��[c���	x'��)�˨\i�հ�=���!M$I.iI���qu��͢����:?B�ͫ�����nt� �ԟ<)��֓�	��(~��.ڿ�^���|ޒL�tmJ��xz�� ^E�� ����zez3!�Sgu�¦4J��Uc��y������cvF��/�_�o|O�kF����)���;��m+9R�I^�Y�Ύ�����~��Q勧�6m'EH����0ޗ���%ن gJ?����<��|���oN2�׭1���cSΥ>fAU�Ϝ��->K�Җ�l��s�~����4�zc�]����o����5������6�Nwqc��a����6�f.P o�E���v�K����{�f�`���*�ϣ7e����Dg��t�]Z�x����ChY�gc�ᶝg��	P+H��p�d�0_��f�ع�k-�H�oŗ_�_�:ʨ���]]��c
Ά���̭d�K�̂(����W�I�d	��*-���W�M¸�޳{�ۊ�3M4j�y
����y�.���\��l��k�i�W�����A��q�BAh芓���.�fq࠰�5�^���0>�F=��5��W���{���ش"s�$*�τ�"�����T�����d8��!������:kW���}��y����ޟ�2�� ,�Ap�[iu4��G`�h�pɨӮ1(!��ф���(�e[��Jx:�H9��Z�U�on����Q��u#O�Y5}���Y�������O|���\xi�2�V�/m�sFg��J��0�8�x(ݾ˶�O��Z�2�oD⽟y��~\Q�}[]�<ݸ�y�8��$���NH?$l���P|�7��U19p���=��)�R��O.��Æ���)��:U���:̨N�g���s��w��!P�o[&Z�Y	V6� �uT6�ϖ�/�p�h"�D�b�q�6t|0ZoG�)H���@�6M�x5eUM�q~X�IrC�J&^���D'w<#q�KZ���1_�ԚMV��{C�3hH��Zޞ�t�>�l�&�x]7ݏL+@@-ɸәt���o���>����O8��PI�B�'	�l~�[ƛ�;6��L�1�,�'y�A�?w)�"���I˟ڑ����f���+Ձރܷ֝}�Ib{u���?��2{��"��7�|�uӡ/B��7������j�z�0����t���9��-�q�}�������i�L��t^^�?���r��zA�7�����&�{����A�RU�nTU%�h����Ϻ�£�Y��̆x{��_R�:!�}\��^�m�ao���ČM��v��<:������i�"�p��	�a��}��`���o�E$�$�T�r=�@�T[Od�ݴ�p/z�����:�1�roMR;Hj8&*���>�/ѹ�`�>��s�X������l����r�@Z�fռ�w9��铮�E=ѥ=�d��}��@U�F���W:5����#���t[���FJ��KKz�/V��}�T�҉PO[��	�A����9B��ղϩ0x�_0Sr����K��!��4Q�jeN���7U4�o��Y��p�a{=��X�AH����"����?�c�4�>�]90Be�͉S �/�-�x����v�eG��wm�f�w�%J4�⟭��Q$��k΍�P�r�CZ���c���L�m3�1�x��9��t��z/�V� �<�/E�3ly�c�F.�?8	b�}P+�B��M��J+R�
�4��6�=(����@�!%e��+ߴ��s��J@���DwIK��Z��0{Ja��[�,��迷��J�'Q��w��g3c�E�1������I+��ϳ%�7�\P��6q�K�ͫo$�R���^Pdi�*kPQ��l>&�c�CB�*�=���c^�J��5��P�\�
E|	����I�L��<��C$ ��!#�qQ+I�&J�C��4;:��,@��[�7"p+?����!�w{�w��<YV����Q[�@��r�	�Co�W�<�*y�ls�M͢�M%Va��
�~}�q��Љ``�7_}?�8h����'�C)�=R���&O�SۊϞ�	?��������2��2~L/ńT�Y�WΌ{�ɸ���eЉ�E\%q�BA���
,�/��3������K�C��*�fv!̛5r�!��D�/�#�QM�2QX��*3�۹���.����;���dP}_ߴ�M���=���@��_���s��}.�u�$MRdH��>A��ndn6���Q�.���)oF9�o8+���K�H2�Mށ/ވ��tL���ť4��W��q~Lf�E��-8i,�0c����
�2�y}� ��$h�d�Wa�����A��7�!9��jW��ڴ �S�g�L�;���05�{�-��X��#��b��+������ ��
�ԂYv@�q>!�3^�@�U�q(K�a��=�e�1r�&yGr��@�5�c6���p�(�
�ll�u�A��8١�[�?�ZA/6�>�5��Ť���f:E/p��RZ�bGe7���0
r���=~C*�-�^�`EH.񼹴T<��#,�"�p�R foR��a7ty�(�*���+Il�¹o�b��S��f�����l���0jا5��\�J�s2t��H�N�(�/�6�h'~�M��x�u�X�j��W���i7\D	h(�+Z5^����Q�rRE��:�p>q+����E\q��0f,��gG��9� &RP����I���p���{�(}�c�H��ˮ�-� P��H���*ж\";�;�[�(wb�S9�F谽"ݷ�A?�hx4��Ҵ���J~,tM�S����$�K
`�F�X�A���B���m��$M&��,�X��sa9!Ǽn�j		QL�ٓ����w��C2��);;;��{&=���2�﵋`�l�F��U�]�pI�!�f.6L�r'��'��Pۃ �%��)z�|"h`j���B5�����h�-�@����6#hF�G��ʄh�5��q�KL΢S2��1�U�Z�.Z��b����X/�2��a�i�M��^��8`��}Uk��Wg��jU#��#�P5k���p�+1�����h�oy5d珕Q��=��*�/��ZOȍ�wr�+�nD_w��-^C���X����r�ٓ�F���a�U���[^�d�0�E���k�n
�p�j�C���Z�Ժ_a�Z�4t��h6�8��6Yl��>7p�S*�p���G���k$3P&DݦT���z��]���Pe8�Z4�xF7�P'�h�`Zͦ�%�|�����T7���:�V�ˁ"%!  ��UHV 9X~���.����MGP$� ���0���B�b�U����8�)3�-��T�^��5j^\�$ݤC��d�T�v�s
I��`?a0�L��:�f�]�*U�j^��̼ ��㞚f�� �#�[��XE����O8Z.�Z��������!p5��+�%3.�Y���gn�����)�q�n��k>�x����/I�
����e�?����+���C-*�������~p~c?Z���
����-|,�Eü����X��7�v�`�t��6]�/��9V��f��܉�l���t�<T+��Ƌ��&Dɂ����ۋb�G�u�
�؎�hNy�:-->�r��9����װ��N�ςZ��	mJ|ޓ��DA~nmy�M�Mre�S[�o�#+���>���W�I�Y�p<������BK�={�cܯ��(��p��v��%0��c�-Ww��C�A�K��X����́�H���X�5ݤ8�<Hѭ��?]{�t���-�p��v�Ł��9��t�V�� �7�(���FlNFC�2�v�QQm�-�f&��ơ��"vJ�=O=�,�9{gx1igJ ���zƠ�)A7H����d��6�R8�����2b�D�
-�?��Q�3�~��&��g;�XΚ8~�a����(�8�Oc�7h��P�p �ˏ�.D`t9mV���V�� ����A�������F˃o6QՃ���	��t��@b�:~�~�CO�_���:Gz����Ď��������郣O���z��c�m��;��z[ ��n�@�B���sܔc���Y���s���JH^�Yy��l��!t���A���jh�j���JQ��vo��ISTR��_7�}�'g\Bu�y��
�fz�!ڪ�2�l1Tg%��wx �'�T�:  �K��'!�^��֌L���H-V�V�_�F�H	(fFtF����8e1D����6��#�&���<�ޥ/��.����X�-���m�l=�e->^n���i�v������f�_ h�����oAr�=�n��|^xK�J	�?XX<�aL�#�5`�(Ƿk��_��Oo�$���6� ��(� �Jź��U�YU�k=��<~�6I!�kvh=���ӥ\eDx$v���]o*/t����ol���.2���@��U�jm�d�!�ϛgվ�mk}���g���<�у ���q�v{�^#���[���3A���u�_|P��U7� (�m&A\J��5��u`+�..�^̕��S�Ӧg�%;*�4܍�:ձ��� Ȕ�8Kђk*ۿ�wD�bF����¼⠀1G/f��Ŵu
�6uU��)�^��+�+τH�5C������� �_l�4"�㸃�6�Q��V�	wqq�i݆�?];��{ +:t�ږJOo�t�ژ֞��>n3�_2^�zF���N@�U+��8��bV�*�A����d=�@�1��;�.̜��f�9Xd�{�*�:��H�Qg�	Az��6��%h@�?�.VB�$���C����1/I�S$�gf�=
Jr�y���ƞZC�n�\}��1ܓ�
��V�*]��m|V��i�.N�nTT��v�W��&@�ƙ��H� �U�P��Ȥ~�褠6O��km�P �Qm��گ����[�� �����l=ʆ�G�ձZe����b�%36��
u��N��{f,ʍxg$Jc+���+u�
Z�2�b�Z����Gǹ���7�)^ ���)�UG�,�_#V̧�5�ȴ
:U�]%DB�v@��`T��n���ǩM�u~�E���ώ!��ǰ���wؾ�@��{�8I����"�Σn�h��G{��8�O#X�,��&J�t��W�����y1�p	�Q�#��ːF?�6�9Ӈ��"�#D����8�Z�Q����]`��n�
/#f}0N����rب�h���R&�fP�$ ��T7��7[7|�:~�dl���)��T��_"�P�sVL|H	K��ٳzX&�0^���M��0�S_�ް櫧�D*��,��1�E���wj��̈́�>�e)<�I�@��B�����L6����wؑ+�љq	�
�2��mQ}/�7$��G�[0��^��~�kW�#�}8�� :�m� =$�߀>-�k�J!_S�#�h,���wh fL���1αx�lXG3������ҹRֹ�>�����u7G�E�e::���o���u���W/�����	��x���ۅыu�(M�TN��3E��q�qϾ��p��6\р���1�}H��*O_Z ��L�5�ڢ�\��ُy}zL��u�1��b�0�I�8;3��D��n��]}��~�7;HΔf���7�*�=U�W�]
����.���錸�d������g~FK��céը2͂�_Ũ��P߸
 (�!����0���>z�|���=��!�XC�k��f0^�ҳ�I�,���`�5�����[��C]�Ab7�L��'x�jYh�����-7�ӛ%r3�9[�!b�N8M�̫�ؒ���r�������i�Mv�.�Sa@z�!�Q*.V"�N���O�Ѩ��} >�gS�H�r>v�����IR�ӎp��q[W�J�R������UYNO�A+� %��eڱ�3@�1���W�Κ�����VJ��(-�����xD���U������ڃ��l��"N�Fb�_MՌ%v�줄fp9=ĺ��;ed9�l��X��}?!�:�p��0�HQ�� v^�K(e���ᇏ�������Ǎ-���x�96������T0�6v��a�&���j��a${�<�4ן��XK��8��+ȴ�܉4� ]�:��ѻ]���}D�z	[iIۂ���sYhUyY�|;fT�@*�Јѣ�օP�]t�M�'��u.(/\�E���A�/���7p�!�����Y�Z#�CM���ue$�b�X�63up=�b�i4��AY�5��|�9�p��6ēsj}6��z��U�,���;F���0Ǹ��C�9�����ioX�휯��E
˳ML�ï_0.�|�/�M�~���@�	��s��Kpd��"B_pk�j�=8" p�:-�$R�@oG@$�ʚ��U�q9��P�  ��~��hlr4do��R����0V��Q�넯��<�85��wl��`����Ɣ��.���7���s��%EG�ȵ�j�G-�><8��ǂ��ˀE��f�}Mx�}�  Yvj���l�t�4�㠸��}P�U�yk���W�G���E� ��y���Hn�׈����BZ���C�`"*���ϝ)iv�D��v(,]Vt�l�)�n�JQDjBwx��_���<�	#H�nWMQ�=w�}$�� ;�,mR����������w�Y<����,��1�*0J�J��H8P�Ը�Bc!�X�#Q�z�@�>}\�%zǟ�'&q&�t:P��q�*�7�ԠS�lV/3��-�%��.P�����C`��t&/4��i�8Q�P�u.e���u�l��q*8S��z�GY��F1�M���$�&�{�����׊~]�!��|��ou�DF�6�eд�����v��R�3{P�:R�����M;��#H���WXKW����x�1Jԉ< ��=���dm��C�2��U-�+����h=:��N��
'�LQ�/	�'-�~� s�ѣ�k��.�N������C-�����4ʞG+!�5گ��1E.�c�:*�"B��#%�4��=jQ��%�A��n�³�c��/������Xm�MPT�CD?Ȁ����A�k��ʑ���.1�"Q#�
�Y��[�.Ɩ�Ո@	�R��2D���R@9�Zy����F2�DA~�,$�6�c3��촟Z�~��
���d��ㄻ�M՛"�?�~�:�w�b"�x(�$�	������K $���7Zϴ�ynP5�.d�����9�E�0O6i<�����GB{s��cqft���:oa�+B&&��>EJ�A��9���p�,p*�0|��?�ƺ��G��04ɝ�nHG��
�ϐ�[<���Ź�I
�U�5D�k��e���!�����#0���f!P��h�U��K�xTo{����_�m���>Y��v��݉��w;U���Aw�Q����@�{@�@��V�[i��=������q�:�Y(FNM +�مq{+7��_��Q�<���-5?Pa��k�hdv����Q��k���|I��6�� ��TƟ���ؠJ����򹊩�@�L�`�������V�G��]"$�	7-lQ�{q?
ZUβm������רu=�PS�%qs5�?BA�մ$f@�Z�Bq☘4)�:)�sK�0ȝx٘�BY����"T�5#��bDe<�f���]�N� _��1�Ed��=�Τme]��ńV7�	�h�z?d_��t�}r}�~�4@�<�i�t�R7u�
�\��]�F��������P�p�a�1y�'	?���W<��ş�qb�H�~Њ+�#��tf����!�+6��8K�����5vG��L��|S���T,�f=��I|L��u��j.��U	&��5ƛĄ���K�][�L��&���p7$o\�Sc��̸��c�o�P��uy��=��4$i��>z�����^��Itv�6�}�ҿ��/ֿ����d��J�Kq�"K���������F��ݪ��$����2�{�q��~�2Q�=~s�o������ r[�ڥ]�q�X�oG���{e�XNn8M��uJ�?�tcyi�v�oO��¹�z���}��ٔ��V���i��0��i����OhE�b2�9����q<wM�d*J��"W�6L������~��AH���V��7d!S��=\]AlO�|ތ��V�-C~������v1tI�g���m�4,�I_*��DЩ��J>�<����v^�x��k;�a�`m��q�~JQ{/��YX�3�����.�d�)�w�y�m�Y�����n{;ץP/[`*�j�e�[dͬ��n߃�P�I�[��J9ل�"4^�Δ�V1a$~�y:�!tل^�+�G}O�����VBઊ1D��6�<��_�rImjα��Z�6�2���s��d����08�� ������Ao3�xv�g�{���R떩��k�H��<���Uc�*�[��G����mF���T���V��HǮ���]���X�Iۧk��,�D,�����2ӫG���x�f' �{���phRF�纎�V�����4ܣ>�����y�e�%~�h�#J�B��w��dd�$0m/����Q�:~d
|I�ꯘ-%��E(r;{�vϼʹUA�����v2�j�%�tdεrVD}�w\�P��m�O̲9��������+l��4O4����).A�O�ʨ2�d�V�����%���)��͔�@�a��W����V���т������O��J���C@���H�GF�ʰ_����X9�����/� ��,�ݲ�28�yڗ���ř�?���������DEsg��N�9M�Y�l&�VD��Cv�K.�Jl��
�Oei���gK���tS웞�I;���a����Qc��M��ҩ���厛&�
�as?�d���	Nd�N�vi�Y�0��A��J
�?\A'��������;26����;���p�tW�f
o�B&��Dɮ���](����J�-7�)�,]&o��*�Vk�o~Ov��+a �o��Q����*I���W�v+��&9xK% l�L@ �c}�E������N�6���L�a?�P���lU�dǵ�52+�΂p��s���s���f�463�,TX�d��;JA�7��:�y��S˪�eJ:�%e�xf~T�s�/�.7��!_L�b��J�1W��P��o}P����NUdd�!]��$T�����ؾ���[Cz�zd�hU��?}K��/�NB��%-���e3��dGcE<�K]բ��Xq�����
�����6_FY戮Vcx���,>eW�PWؿ���/٫�Vה~�7&ܶ��Y�����~}���v=[4љ��Qe�I����x!��%QU$zaO_ᢉN}�;��2��o�����Gb+N�ͬj�����hM*]�$|�T4��l���X5
r����
ul[!�wr��G�e3��9JqI�&/�@Ǎ��U�Pp��7�3���n��O�Oy�;A�2yb�ؙȚ��� 2��P+/
�L��j���6-����g�QR�����9l=��v o&;�.6�I.�����8��%OB5$��̸ה����s��&�D��bK��$S���ׅI�|�$9��gZ��T#�MC�]�TV;�s��L�2��&j���3�*��%+�
��{�9
�$R� e�p��6�m����,V&9I
,����A�Uw�i��3��Ǚ<�,��C��eoۼ����&����7������c[?l���;�Y���5�-�2�d�'H�z�Y8a�j�)�ЧE��4���(Y�/`p��L�/ۿ߰���|�f�̉�o�ެ���h�8n������*+��`��F
���
��k�S��̪.���O<�-�j4��틚�Bݵ�Z����������D��1�݊��ZU�Vz�)���3}ie̵����Gu�,V�g��:�5s`fE�B$4�^�7� ���<W�9

����?�X*�nAd�W4��l(Qb���Slv�\�G&����D�'�a��d>Ɋ	@���q���X"}��$�π��]#]�i�ifK��zC�jQ�j����/�}��:f�(������Ѱ���4��Fi���n�đzb�H�GN]�fu���~6^�=*�dql`m�N!���ѾS鄓��y��!jՆ��Y�tg�Ս���0�y1�H-g�da<�j�ڵK�0�}CdόH�C6
��8��e���l[�[��%�x���k�a%�7�R*�4�(VaO�x	*y�S#��Jʄ����d'��V�{��} ��%��zRcp ��K��fN~�nҏ�4yPRU#)�4��+�X�ȉ��u���� �v��e�H�i@@�ߋR)�h�a�(���,�T�� h��2��?L"g����y�)8�������� �"2�ae���?Fr0�Mg��:���@K_c�-���x���1�+���>�Y��x���a��R�<��(��>�r!I�������R�m۶i*K 1];�S�z`�A�8�#-!��3�A�I .΅�"hp4"�q��=;|�ˎ��0������~c�|�JAǂ{��+��_E�S���0��c:b�V��1SN>��|rKs%Բ�'A��ۅ��Gsa���u��$S��Q,c��(�o{ �ɺ���������.d�kR�J�&�* <�W֬]�+I�T�Y�e:�N��6Lą����49� �7�t���J;���I�6H2��x�
���l٢yG ���q�NpEf5`�ܑ���p��\ԈfYKm�93�p��Y	��[��V� �0���A�i,�<l�
��C�j�bH���D;ܘ:�h�ΔL��4�������������c�DQ��	q�r�~s�a�<��%�Mo�\آ�7r�,\��;��cTǅ�1��;'�oN��%>�N�dOl6S����8]KN�SsS]-)���i��?����SH"�#X"�Ѩ�#F놲|����4�Zo2.JW�����SU�Q�*�
(/ѿO�e���Zo����X���C������?�����,�d����N�����Brx 0���&�s�� �6lP����5XU�"bsu�	��Hb��T�qR7)QT2�pT<8��Wi�`��������Y�eX,bڡ�x�k_����.���j쏥������yC��]� �u��cB��P�z�pH^�j��?�fy�:y�O}Ɯ�,����D��G�AlݺE6�y�a�k�I;&���-n��<$���+�V��ɌVӕqN�Ľ��%*��W�xq¼�H��O~_��H�
�C���[eϋ(1�0��eX�[��+��qҭ \m�һd���i�݋�a�~l�TO��o�,U���~�µW�8V�� �}�k�����`mJ/�㔪P|�����Pc �.��'f0�0���Pc�҈��l�����0G]
���|��s���8�%?�D�
���ZY"q�h�0ox���V۲ap 0J]#y�\����Z�!�g��i�J�u+��f�������xg,1�אѡR*�Jo���3f@�W�W`:o�T���?W����]2<tD
�b��j�>��P���XW�f0P3?����f9n�9�d�n	��9X��K����s�>��7� _� H�նo�A3���yC|y����Γf貔���19|��3�ʥ���A�b��.��K.Q�
5�����Z����K�@LLw�xu�ʀQPa��ΦƤ�b;�(�3�_y�zl\�#S�� �h�'�ö׋��nh|�%	�	�7Ζl8[gB�da>�.t=hVN@ðq�/����P��-oy��p�z��䤑M�n�lT��E���n�]�xܑ/<CN[{�T�jR�c�2&=�>	¢�A��w���$g8����^��hr9�%��#��NH�qQft��.��Z��J�]��ǂ�<Os^pS}p¾]g���s���]ق��Aw�]�Y��5	#�T��_��������37](=}+e���%�sE��Di��D����*���7�Q���p�
��&�^�O�N&f�>q k�@�Ŵ  vu���0��ׅ���،�f|��ya��R�to81�
����v^0g;���1�`���K����R��
2b�ep����s}���	�~pTc@lc�Y��KSy2:,���o�CG�w\w�|��~P���Uw�-[P��S0��]m�!�/j`�����5�r�I��(@�����c���5'����QvfLD��ᩤ	�%��6��d��~>��d��Ȁe;�f�
	WW���b�D(�Ұ�;�U�����|�w�I^}�:�$n���:2��1B�';T����'� ��xF��o|C3�x���cB�L��+-���4�j3^���s�9G���.�/񼸨n�q%3љW.xիe�V���͢��Au ��2�=�VFZ=q�`�X*@O�

�y�# �����1��� �=�EB�C��&�r�3v�z�/ˮÆ�#׾��r�Ƴ�H�\�=�R�%����*�&�M7��?�>�cϑ��X�~!��Z�Ɯ���L�)�SK�|��3��ɖ�4�C����$66PR��(�hE��|*��'�#C��� ��������o���$\Q���B�%m�F�9X�|�f��gT�|vK"F}0� ���C���j�ꆁ�Z dۥUki���QË��0 j+ �m�]gc����0�#D��GG�sww�,�]jf?T.}	����&�B#��J�̐K6&����� U4uv��^`� o4�u�E)(��`QEóL	�aG�Ql�j�բ�9G]�
�ɞ���W�R(��q�v�0`s^YC>���F(�rA�"��Ss��2�R3$���F��o�'ʼ�� ���V�?��@��/��� I��]� \N�1*���֌����<E=�4�����_)Fz��PS�����N8r�5o��V����~����2��GU`�����) _���f׈㱁'�_i�L��k�E�8p>X�~�NJ4��ڌ4�m������zG@�~\r<m$���u��S�݆	�c��ƺ񼯶���C���vyp��1C�AXN��6=�e�#H�9n���`��=�Z <���F��$U���h���իW�c��_UU\x��rҼÚ3*'��4��1���m��ҩ>�^I��7�Y��̘�4OE��(�N_+�����^Q���,�*�d���:>��
⌗%S�5�A'�|4��+��B��?���`��ַ�>���W�E��:^ ,Vʬ����	3���������ň�^���o�G�Ŏ�B�2Ci��P�HB�CC�T�uȆP��#�^�3o������6"�p\g^,;`�c��g��n���m�Ш,�d�-f�p�GI�RW�}Ǖr��uf�#f�n$���<z9�!mCL.���%�񔵬BC[OOY�v��r�]�I�5�4&�=��i�3#`�
�&|V*�R5P����w�m��,�l4H���"�5l�>�� p�+b�R�����a�TI���+gd��{�n�u;Y7�0xtl�f�p�+�&�rF����l���0�lR�,�	І \�6��a	�G����+2�z-��5E�Y��=��i�z�5[^�.Eؾo�R�a)[�H,訙�r}o./s�mFiƒV$B.�J�,�l�X>�W!�����w�������a�:�I�/pF{���p��+u ߫��Zə���L��u�8�]��.�i{Eثvb�]�3��ZT�;n��av��f�d�t�޽gwa&r��s��!60c����KVb��	t>X�}��j��1z�3�ZSt9a�8�l0�x���L��k�&kVwK�ё�ډF���U��w�j v��\rɅv��h]B��a��H&���W�z�&9p�jƴ!l^��ƀk�*X@�c�Ft�}Y-dpI�� �|���U�7���M]/�����`a%�&��z`K�P�.��L��8�N^!6�0c�ho���%/�̉�����C�>�3o�G6k3P���8#��f�t	ܴ��Q��.�@����/�J�;�S�>h�d�Ri�hJV7��Oh�=/Ԥ�1�kʂ0��D��U�ȴk�I.��,6���!���c0�oɀǲk�a�f|�1y(�+A\��K�Ы9�%�&Ԣ�H8dU�v?�3�~��o���b#F(1�0���hP&�5p�2���`/�ʳ�C�'T�����̰�l�A��۱=NB�"�v��.v��e���
ɰb�e8�<�����m	�m�C�d�� t�p��<%�����;��N?��׿��e$62�����3�f�.�8�!��;����Zal��e��r���xE�D����9�����$���1|ė={�����ʿ��0@\It�KVʅ��L6l�,�jA��T��	�1�`E�m�ZWo+�(`��#�ZU�(�*#�@����/�O�Se� k����A= �
B�0�wbڝ�{L�>�1��X�Cg����Q丵�/�Ӥ=H���i7|�Sdͩ����v�B������22[l�9TS4
|�q��)�/lU�*h�x@sV����W=0ddT�R�����k*g7;zNϡ�2�z���{�,)���dd�%ʽ[oאK�)�z�Itù��r��a�a�xH8f:8jخY����1g�UW��zVv�8"Q �.Þ_H��bdT��.��	CM� � 緼�M�w�K1��f`�ƍ��g�����4M.��{�,@*D�­1��< )	&���`b���1���]
ޭ�֧%S�@�q���5�46<�����Q�W���iz>���'b�`���@��D�!��@��Q n���xȀ��׽N�?�|M������w�yg�˂�Y>L>�l_G�(P��Ǝ�&~�	{w�'G[��I%Yg����r��bѩH���c#����#��`��}��zV��L`G�B�a��ˠ��/�\1*	�{�W0䫮z�zI ����؏!�XM�}�ٺ��k�y��3]Ѩ"a� �
j�B�rg$�Ŗ�����W���a&�)Kr��ae�o��W4�-"�1h0�0���m�f��@( �3�T���x���q,Ap|���~�#�aψ£��A6��j�v������M1�tH��}�谖zA� ��A��9 ~�J��\��j"����� "߬$R,��f�r�[����%W	Md ��{����1z��3�Q<A���J� �
 @�E�[F�# �XK��X���Z�� j�0#Ѓ j�'Ӌ�4�[�*�xܡ��ry��u�}����I�q�K��0U�/]>(��|��iш�1��64*��P�c{�xA�ш�1�ne���́m�5�|���Z��m�{��#���Tmd\JT'C��K_#KJ����J�����{�O?�9��iL�	�{G�KS�	M���e=����͐�-j�� h�#�[jcCK�s�Ӵ�fm>�I�'���'O�'*K0h؞zz���茡� ��ؙiob p� `#	��h̳�d��c�j,�+o�\R0��EѬ�x��	 CK�(A&qs7�x����4�%t/�@4
@I��x��2�)l6����l��m�+N���ַ�_��_u6�;�� �i����m<���MA�v�5]��W֟�/���R�nؿ����zc�lT���@��K./S�ll1jۙղ?"�#��ϕ��/5�-�Zݗ�%�dhDd�Hu����%Mx�[(��N�8�˞k@ژl�bF�Q��>�W��W�{���El!#F�3�[L� !�*$�O`â������r�2%������)���Z��n����Q�)4 �?�p�P5п��@���ҵ��I�[�:�K�3-S�Q���I�c��M�����5������w�*�x�2��WF��(��1;ʄ
��
"�\�B*�]�t9R�*pT<�R��0��g��R.��z�e��f�4��Be<	�e��Z��|�{���!���R�� G��2P��f5�[n�E-��#�T����nE"��(��W�?2d�A[S��xއD�Rr���& L�\�ׅՑمpcL���7�$P%@����K�.�m�&�=C������N�n�mG�	������n����\�����~�=I�;�&Œ+a�O?�t;izG���\���}�q��D����O��/ɑ��a���/�B)$KZ����a��1�RK���$�$\d��![�1o�!h� �Pi[X/��+j�t�������F���4@8����Փ��F��t�F��(�=�ܣ���p�`��t�t�̺q���g�Zb�b�v���
�\��������O�o�2y�������T^Օr���Q��� ���AF8�2�`¹�R��x��Ы:�P��ȑ1�η(O?�O�9o��
��QU�Y�J	p��G�3)����%I��	!���{�fDw�$�D�	�� -A�o&i��JX�]԰-s���m��(��t�����#L����F�����Ibv�#��IC'�r&�a�N�v @B�wG�@;����'& 3���3�����y[���;�1�Z=���4T���!����3��G���p��cN+�%�s���(��
�� %@HT߈Q�H��=���o�A�8��B�*w�X-�4��G�=�EŜ[�h����e&ۡ'�"@�`l7��x��A�q��-�o��D���t��'�5�ˊ��VR�l$	��P�	�	�V;C~z��4�����!�M'^����%S^��G�=�xiE�$e+�:Z�\���hM��ukd��^��	�F2+k�'4:��xE�"���\G��	-�M����)yAM���a)���c>{�OFd����_��F1��;�D��h�U�H�^I��m�I��u,��b�h<���`��,��[ u�+�x;���ΤF�i��m~�#�:,ms7�RLg���Sh=���Ͳ�6�O�lp���.�ț��Z9}�Js�5e�����ۼVPȓF��rѺt,����%cY�r���(w�����0���+H���t����a�Q�
ؖV�7������*�e���k8���m�4 ��m����i'������
Ϳy�������W_$�>_F���oH�kn�%%Y�AA]��¹��2]7K��g����Uv|�����V�%�Ε�����=�<%�m0+��`<�KO�Ig�
�)h�iE�:I�l�j�6���,�-��`ʻmwޅ`��9����Y���r�\w�I{���kd`�82:�G�{��F@Å�HZ��UU��Ē�ͽ$ryy�L�B��s�(��q�h.n��W�s��^s� w�X���a�}�[8����
3�b!d*�k�UO�U��pڗ�H@p�}@a���YҨ��&���hp4/tɮ���ޗ�S��}���+�'}��_;��b�X�#inkʼs���*���o�`�R���3$�>�TʮV$�`��nCnP��W�zz*j�����X,5UIƴ��I:n���$��L��|�$l��C���eɁ&U�hؤ/?���Q� ��G�J��%w��7f����J϶ *�\r9f��T��������/_�Ï"��z�R����.����H�>f��"�_xN0G�1\ՌN�Jq>e:㺵Js���)��Ubs�l!@��jvA>Ɔ#���5�����ȣ�J����+���74K�����D',	�p'�c8�8'¹��2�N؝��Xj���Q��P��[��CU9rpL#��9u�iV�������Q-�nV��Ɛ�m ��u[U���e��j'��Pf���L8.��G=��[�k�B��;�=�Tn.s]6W�G��U���=*cպ��`44ܐr�Wg�(4������)��șq./_It��JQr�a�%�u�ZS��4�;�P� v����n� �u;�-��خ��v�9[��h�ߵ��>w�I��LY�PD��$�,l$��+4��&J�-�I��pa���Q&L�l�윞�R��J����2:��˨��<�s2u��C��X�A����eI��3�_�¥c�Xv��oZ�dfq��S��d�K�z	Cfs.����
^B�ό���O�r14���{��J�Ud����s�շ��a�F�s&c�d)C�u�L�Ê��b�[&�aUb k�� ˀ.������z킟�1�EG�d��$���a��1{zz�Z}̀n =�.xhHZϭ�՜�ņFBR�(~G�
�Ff8�^D
��l��j�T;п��!8/R�m۶��}�X͆-� �cr�%�ȩ+��/c�vH
^Yv??,���#AL�k'�aU�\���[�	���<(x���m���_s����(�����JWπ����@���$w�nB����Gi����d���$��l Z�s3�Ta�c��8����-xEl���W���6�+�0�u��o1��3a���&��PNA�4\���(�(�2�#�rc�b�ID�����d(�<�c,�^���L��kց�I}���=��v�{v��Y�j�,]f�����e���X�W�è���!륯p���2�U\�9Qn�w͊�e��+e��k��2#��,�{�"8�l� �w<I�kV���s�	��I�ƒ��E6��DJ\֤c}8V� p�եy�H��w(���cH��c��"��� =/����$?�b'���E;˄����:�:�r����~
h�,�����9���N�c�[�7��;��s�g����Td3_;��L�3����s;>,6 ��m��dQ1�����|�;?�姊\y�y�Uꑣ���<ui�m�M������Aƽ%�s��\���
�7 ����i��C>b��3r�+6��ҵZ�hp`�2������Wj��昧j�Ł��^�n���oЂ�x������T�A�3���F�!���r�RG^x���e�&� �ׯ_/7n�ԙO<��w�}
�L��4���0���.��eH?WR����ޛ[z����Y�K�}E��,�UHB�Y�&���ej��$q2���d<N��$�q9�	�+�8,�)��n��lV�f�EK��u���Ϲ����{���,��=}�{��Y����w�+��x1�����ԧ>�0av:���ݽ�,(=̗]��{�2�=I�u�<��:9��9dÂ2�d�����`�u	|F��]�I������ҭ�}N�շ�b�W�SZ �����56PE-�k<L�n?ŭ����LZ<:H�ƽ����|��7��[���q3����t�g���n:vl13�L�23^�2��U�y[�l��:�x�С��]Ď
̴w����Jԃ	�b��|!��`1��Lވ=���ݟ��g�b�A���1�y��:��p�ȌwRQC�; ���W_�����%5��vJ�U/� Tt `L�|�/{���������Ed�2Z�������M8�ߙ�]q�tF�s�F��4�ޕn�w)���>�^�ꗦ=yw�͢�5҄�6ƻ^1F��~������=>6���o���{aW�0:rd9}�K��y4��}n:�A��Uu���@�Y�0�5��0w�za ���//�-�+l5�ھ��o-Y}-��|�W8R8C\��XU�n8U�w�W b�
��`Zވ��q��B�TuG��d�3���b�W\�b�B'���Zn�����+��F��1�bԀ#�]�a�9�
�dԏ�D��3ϝ�nF�#��i���Ӓ��V�6G����#���=�Kg��V���r5t�u�J��ԛۮ���%������u�f6"��jf��↶��F����%(������{~nO"���)������!zW�L)���^��������Zv�.Y�^ı�_�����fS�hZ]j�=צ
�R��O}j�'~_�3��ߜ&�\cm�
 .���.�����P`[r^ r��{��ǘ/�݉�s�}hV�P���k�413:">�q��Lci�%[�	O�y`�=x`!�����w�tɥ�(;�m?��T�^�P]5��_i���"��On���V���[�A:ppoY(`��$���bj�T�r����`�a,�{�����׿>�����9sPi~��/�(��z`p@�<N�9F�� �O�g �#<ª��ک�� �:a�Ӛ,hְ�o~�bE���������Y ZU�_��إxO)w/��ӹ7�x�D�s�e��7��嚟��g� V'lֵ뷊� ��j��28�<7;H��ޖ�>��~�^�'P?�:�i�5̬??�p!��$�ο͢S�-K.��1���[�Sth\��}����y4@F?m��ڧz��rQ���vjYԪԹ�"vI��F��4�8��L7-�׿���;��a������j���4�5J����Mb h�8�=I�UJ�ˆ��R�N�Yi��S�?%D���h3��*N~��wx_�)p��7��#��qb�y�0����T�h'l9 �w} :���x4�-�-�8�-��~����78DQ�?�y�+�Cf�!�}�����ɶ�K��H���_������M/y�3�����_�UE��'C�U#�;���m.ޗ^"�lKL��;n�N�h���X�Dd�n������T��g����\��Y?�T5~B��������矕�ߟ��|� EY�̆���I>p�#�-O�w���~����{�-	�N9C�DL?ap�ȹ�Pe�u T�j'�JǞ]�I |�q�� VQ��j�Ӣ��6[#
����J�{��Ep����=g � K�U��P������b{�7�]��r]�Q�����¹0���������ƸX�^�i*��p9��k^�Ͻ7ʹ3+~�<8{R#��=��H�J"�VI�<U���$b��[d��h=K44r���T�	&��]<z�ȸ������v�"������n�yN6Rg���؎��/��@3-.U���>Et�ra����*��!w�|�+�}�J	 }��^W�v�3k�H���Z*�b<� ��wU1�.�<&�%�h���[ �ƹ  �����������[�R���� ޣ> ���}���RA���*2�XE���y���<�$��KGsM ��y��P:��a7b `ٺ�hԏ/zD�VTX�,��XZ^z ���I���X������{�M�Z�8o ���/"ب(&��bM��m�yy.&o6'�);�`����[�IVϹ�eO�ux�=�N�� &��4���L����a/}�ۇ
�Y\^���@"�e�f�\�>V�N��M|u-Q���i<#����+��+��ha� 3��,�b�DW�6d�u�yX�ϫ�W4*y�5br0>7�x%�Vq���ye�~{�l��t�ܗ!|�H�´���d\��bu=�N����C��DM!0�.���v$�Gv籜���ă����u_��O�E:�A��]�b�L>W�@{�(r$��%Q� %jy��K�V��ʸ����E]�j�0T5�*��=M5����I����C��Oг�Qi��Y�}���p��jYXN]j�5g�����@��}��<�������ԧ��g��IOf���	�B��B� ��x	s� >��a����// Ѹ��_��_M��dòZ�$K�i���un�cP��u�߰^ū`��5��'-�@�a#:%G�ca����]E}���g�C���9�������i����.�@�f�
��`��ǃ�q�tǝG������ئR@+���#�	��E��䩨� ����ϝ%��z������"Fa�EdZ���u�ұa��i�}��Q��jUE�#n�ކ��M���`���@:� �Ġ����N_���Ro8�v��W���Z�J��5�m٩�8!�vQ?j8CB�s��$aF�I81V!��=���ʈ�bU�-%�9SU��t�[2a���1��;�t�X��JS��aEݬ��q���*������s?�sE����u����I7L��9 !�z���q�U�5h��ǎ.�ߙ�T(�D,/̏4d�͉��N5U'�!�
�'篛�����T9�хq� 6�kâ�@A����n��i���zl5W�ˣ�l:�o���}�53�f��i��+u{��U%s0 ���s}����%����__t�	� ^��/�B���K_��d=�*+s�|1߃8��*=u2�zL�w����T	�����fba~��0&x��߰LK ���/ܴ"1/:��A;Oe9a�Oy�Sʵ�h�r8\�{BC�=G����c�V���y9;w_a���ZNS��}[IeY�n35ơ��;�!a߸Kc������x={_3<�Z���?��	�vr!��>��p;�&s��0�ۿ�_��0��]��G{i���+���t�y&\������'�u-�p�*6a�Q?|�_,ċ(]���[��������19�	Ŕ4M,溚V�^���o�h͆���j��R�#3wX����������V�\X�5�!��%�_��&��:��"2��`��À�d�X75��XIaȷ�r�:�4�2p:�n�����b��G�s�:����k�]�9������/�M:t?.xc_�̊[�,�dq�2�<=����L�i����y��18�tD#��_c��Q� QU$kv����Ltth�5.zi�&��w��=�L��6S���XF�@���a�xhu���UWѥ��t���$}������w6��ką��&k"\7�֫�G����R[�w�1|ٙ��xo��g��y��c
� �|��a<�V~W��.~���RZ��I׿�����D������kj_:t�r���嵚�d!���R&;�ɜ0��}��������da�>D�џ����xЪ���b�c."	j�S"�?d̮9��\�:΃m��a��i��= �k�
h?��9�Fg�ܕO(:��sh����u��Iv��`���>|���$�G'� �)�n�p��x��_]������c_����{
�}֞�g�{ݖ��]�Ϧ�G�������q�S&:��V)-]�p|��8X�N& �7T��G����*0���,��~LT�i��B�A}����P�'i�L�{=>TU�QF�`��p�İ�hP@���gU/���	N����9�*MP�|���Q�V/��-���;�s��ϣ���B6E���e���ܳ)5����s�-H��<����@#�qv�H��;3Y�휛n�클w��|?���᠚�s��
��b_��hyȚ}e�-9�����8��:"��+[UltWaɟ����٫S�
��0r�1���c��K�诺�:b0(;(*�Fw5��3������Lam_��m���{'l��N+�M�/
 �VIgG�'�k��==' ��Qrq���:�I�Ȼ���=�%�N/}�uU&���|�_|�+�
�K�V�\���aqY��|���	�eE���=�š�Ɂ|�^���|�P�[6����~ٲ#:c�����S�]�)�9�ދL32Q�aLQ�u����q�J��#�T�yd�V_�Y�z�D�d?:�K.<w��7,A<J~e�5ת��kՃ�di� ��IdA?�d�3Οh�	� �5�'��1�W��x�H��習���;��u^c��kj!�3c��0����qǹޜ�(j4�o<�)
xUn.���д��է}�[[,%%�$��F����cc�N��a\H��^͋��΢��b�˼�E�/��n�_��0��.�@B�I�p.�n�ݜs�M硎` `����?��q�9�~��	 ��3�w��?������w|/���ki�����x�̍˸���p�*�{@�G�υ(D?�@�L��������6�}d�ѵOp��h��Ah�4Y�b~+7(��5Cb���	�Q�$0{?.n��D�n����5Q̶��'?���JUo�%���M�׍ȹ%<�����_�ӯ.��q������� nbq#s�� 7A��im�0[4r���Gy�U�����O}6����p��x�cӹ�<�����d����_�&m>_�SЇ��<�����@U'@�o�1@���ߙ�V���{^�_ԅ`��h�h�9U�bK��r��
��Ro�Q����93]����	(?���"�
]���O �u��7�u�v�s�5��l&9�'���an�=�9E���6l�Gü Wf�L�t�Э�ܜ^��Wd����n��(�bW-3qq���l4� �lP�0h2w�v�;��0�3گ�GH�=/}���t#�n8NP�;>cK�^9�qa�Ff�y��
�W��2�"G�vL;% �G��q�,�MH��8u�)����5"��ܜ<FՖ��(mE�瀯h0�*/��>c�37P����p^���OfU$l���Yn�;����,U�;��̀��S��?���L���� �H�3{��oHވ̀��Zq�g&ܠI"�wr6��C�;�L i.�p��Z�7S�!�W�}�1�Ҝ(�ɑFh4�K�Q���Ǆ�����ԙ�&ʰ�ȳ�FH�������9(�n4��X����R����\�1H�΄��Q���
 �~���0,7B��$N�i�w�f�4�.��QZY��zG��G�^���Q	Ψ�q%jn���ˮ����7�'�('��G?g�&��)�9�A
pH �}��|0�H�'Rt��.:���rl�L6&㤟�`6���`4�����S}�s�0>��0|��F7�� �|�����I�B��'HMH��ؐd�qSQ�%{�) C@���Z.���/�'j07�>ᚑ�sN�ec^k�+�����=��}�	r��n��e%�Fȋg�3���X���^��X��T��d���֓m�R�;@������R�mi~�=Q!��.�t����VW�\�j7��h�q#a���H+lB?#�b��ߌɾ�O$k )�1`��r3�|�K�.k�����i���=��	�pY��qb��Z$7��}�U?_��xy��ޛӏ��C'`���V^���O��ѿ��22u�V\U��.�-�.5���#�o��]�1?��47ߩvw\�y@�����]|K��Z�Zd�47��X#��%�3��cq�|8�`��=��b���5�y=@�	���sr=�'��1n&61�}��pO^܇@��`� ��K��T�6�,����*�(F��l�8�RB,�8��3D��碿8 ���>�*��d!r� Td��C�ٍ����FgF=;cʼ�xv��k�q�A�����Z��@|]��+7����^釾aL7�i����y���u�hlr|��V\c�H�ֵh�%�0������-_�tZ^9��W�TV�Ro��O%-�Š2�>��������L�N���$b�c�}�ܠ����\��܏���S棛�7��������4���Ä�P{ǖ]v,B��8=3��;@�A1؉�Z���� 8<��� L�2��������X��L�]�RGk�ĐBrZL�ѱt���k_���o?U<�٬�y�\|���xK����c��+�s��Y 0A<;;����d�y�(3��Ȩ��::`�o�0��bԡ�W'Ɏ�(e�dt�������E��Z�z ��4��� � '9�x�\�  	�`��Y����8��XO�7��H�ȸ7�ɴ� ��/�ʋq�1�[�+�2^�J�^\����Fk�Uf)���z�2q>4�,�v���M�f�,}�Z�J����l&|��������D���jc�(���u���^���7�Iǎ�*n��3.4Y�_cCl��h�`�C�����9��l|�w���*PؠKQ�<2n�ĺ��2/�|�Ӏ���uPI4OGe|�h\�����a��Cgk}&�{x ��i@Y���q~ݓ\�.VZd/��5�e�F �<��n�X�巼8]x������4���.�;+7"sX��D#���a��g�0� ��A �=@�Ŀyo Qt�t�@�
:��d<����u�q�0q����@�_���7@������)++��α�ȸ��m��c��
��: 'ǨnBtw�	�	�@̧Ap]�	аy���>�=�T��{�ч,n���o,Z��A
r�`�m�9�
�G�c��&2�ڜ�{��$����w6#E�`4P�M��J-�M���dW��#1���m��7��1F7S	W��O�Of��
4�:�t��OM���_������ݗ�^N�),���3�ɿM�յD8�$9Gy�����$��x�zt���s�����%��8�W�	c�ԤD�9"f�~��eW9�v���'��ڤ1�&�L��Jv��]}��.R��04���N� �N�\����H��ufK3��dYJGg �<#�kp0�1u�<��[�d��hX1����So̱.>����j� ñ���KF��FR-� � E�n:>���cf�WU-<L1\�~���Y ���L AF
�D77�Q��T8��D��F]8��Y@�X� �̒��&�Qm{���g�"�2H��	�P��Fù ^���D#z谈�
��G>�w>3/�~���s��K編 G�����������@�7� :�W��Fǎg	e����=��I��{Rz�eOI��q8�%(� ���u3��z�5{�@jڏ<���{�n*V��Q�F��-~�M�괂���r�Y_E�����;���71Z���X��7ͤ�c�<yVґ{o/,xi�P�`wםKiϮ����V��-�T|�["�.�BTsL��04&��� ��,� Xu���H��Tt�R'U^[�'���ٟq�k��ا �WG���ʱ��\�c`|����s��Z�Z�#(��k��Gi�DyY$ �U34[=�Ϡ�@����ʽ�QﮇC]�eC%�􍢪9@3�2 $�����k���`7�=)��F�8+��-�:D7P6DI���0�w��\^s3�3qٗ�{9}�����9���RI����!=���46SoP�0X�������h�٪m���X����<Y�:U���	��E��J���^w�W���xF7��4�I􈀙�K���.>�.��|��t�m��UG�u��ؗ~x0FB5*�Y�k�=K]Ɩ����+�5	\,,,�	���{f� \FE7����䥩/s#�ݱ��q�����
U�?�������q������ת\x&�	��S]��e�����P�%����iaG��Ёj(� #�� r#]Ԝ���mi����2���ߨO���@�uݬ K%#��|����W\1�ce�@�õ5������_�}���;679U{���k�ԯ3sԞ��J?����P�;�+���l6ͥ��=�Oyj:�����-�O�Ae������Q�3��~��\��8Y�\��hC�<R���g#p>m�9��6��Uҝֺ]*�������؅, ;�X��3Gv��r�{���ߕ��⢴�'k���8�5>n̂U��kTV��+�0W�A+J+*��M[ɱ,,U�|����vk���;�"��C���T�D��!@ �y�� 2T��H�� J�h��J0�����Q�j?*N�o��c`��b� �1�9�}��9@��M��{�e�</��Xm����,un���x��Ϸ�0��o�v�zэ���=R��� ��g>c��yO�rO܃���+����mie�xu3��ՙKwޅ��0�u�iiq%s�,��D��_M_��;���O��*�Oou9u�k�ݴUD����<��u+6IQ}�D�9n�_�P����V�Ś_��q*t�悎�Q[�f��j�	�R�ޏ��Z9���n�ñ��ư��2���x���ΕdR2��;�LD����H���}I��E	u��'lN ���Ɇ]��O5@�0Ѓ{U���q�����p��waEi)�J�� ��|n�7i�.�2{p֪���N���e���Pk �|&+���>��g}J�����oA�<ԧs�z�"�s���_�{g1���G~ �㬑Q��:�is�TZYi�@�k2��H��k�lg>=p�p�x�ymeIs�f����q뭩H�7S�P��dY��{^/�;&1�cں;�6<�>�j���CٱQ�w�����hQt�܈��)z��]���w�?�>��v���ۊM���͋t�'}����ˮT��UڞQ�r��\@,���F��K�]��_�{ݗ�C������{�u��g��M��GР}m#�	���c�e�@�H��]XV� �Ȟ�q�Y�C�X]4��n�V���F���7���]m6*���ٜ 4@��ͣ
�ee��*[�?���+vC�9�q�T��=��<�c�}Y�����97� �q����g��8�\�f��'�u��%B�7���AZ�k璟ɛ,��a�V&��iqeX<%�>;o��"�s
��5Ɖ��/nt�s�"^�}�@=��u����I�N��Vmk�Q�7�r6��Q_Y7Z�p�e�N��q���Rv\�?J�P��ꫯH�w5��0ͤo�ݽ����+--c��)���l1QRe�{���X,�7%I&&��hp�K�j�c�O �jl
?�:���M�P�F+�6Lӭ�H"��d�|�ƌV�D�@8q,L̠��	ȹ��Y�d���� 2���Or��{�J�O�HI��
2Ґ��q�:�ܜCC����;�99��bf�������a����>�zƠ�յN��^.1/�sϡ��q/2f����y��o����d2��F�w͑�}%�⫟�^�����\� ����F8+�uj��ހM4K���q�8#Q�g��W���؅A��&���}��(���	��)u� <�'Yv�F{,���+���޴U֣�L�"���Ț�nRu?��8��1�W]�_WV�r4O�t�y{Sp$�u���{:s�U�fv��"Q����Y�k��i��gq#�i��j
<7� zpO�v}!c�W�u��b�w@s��Ⓟ�j&Q�xt��h����LQ>NJ~g�f܀��70<�w��ƨ�t��i�y(�4�Ѧ��c���{NXolO�1X$����iج�5��|��i�IT�9��3�a�ul�;��^ �^ݸ.���q�D��g��v �����!Qo���XIg�1����J����=���'�o#ϫQZ<�(�`��crS��~�n�]�~oJy��<�u��@c�*?U��,�����.�{��%Ap�E}��w�G3�^�1 �{����w;��0���F���#��ZlG���zb�]`u�v���2>]��M�ڠ����{��(�w�Bz��.K�����Ky?�J�'��+k F���*߽U
Q@@0S��ϲ�Q<e�I-�ɈQ�b�f�p���Km����n@5`�-�u"�J}��o�i�z�&���N�E°�wu�����7cqu2�9N��bۮ�9��4:�ˢ�k}�5��G�l�C�ޓ��M�����Q�yZ��G��j*��T���&��������:P�p�W�e��m�=��m'&x���.^Y��6�����:��e n5�A�hI=�və��	�Չg&"y�v��w�F~;�,��h�(6hx�^W?΍�]Ռ�O�G�VW�Lo��^�~��^��ҽk�;R��0��󰪶<����/���K.�l4�ϚU�{dN���k����0����������2�4���߭�[\ [o���������A���e�ݴ�nv���u�'�L��5�	�H���l��¥�L#��|�ӟO��ޑ��I���/K�?[ x~>��X&@�����	�/�wd���h<��� �$��c����mc�e/��ؤ�9�!"��6a�m�j��G��(�ɮG���&vH��d���F����n����=��\tx2>E�1�ц�H��L��ٕ�{)}�c�~��ǧ'�����xHL���y. b���,�Z*�4����]��x��x�C쿸����"����xYr<W��~Rډ��F`u� 6��nv���Zu�����F`_�~��6z��4��U�l���0?��>����wI��L�=�?;�R�#HPe%]7Қ7Ud���X���J�UPۊFN�EI3�����|����͙m��{)�C;:�̄��l��`[c ��y��C?5�;{�7 �X�aS�?�u�և�
02߭�u=My�0a/�N���O1�x�:`AM��s�Y��W�����7�M�K�4�!�CO?Uي�ͱKZ0Ѝ6WG��U��F�G���
S毕�}���$�ƈ��KM}q���!=���=��6E��g������`i[�ش{8Q�?۩0�킿�4ͮm#��4��ζaq�Dm7$��Q��������3/�n�B'Kγ��[J=Ԙ���iϢ���\�+�*��Y�u�F��f�+mp����_�fTc��*��k�������;�AC�`X�,�kT)�V�Ki�W�^v٣J�E:�/���N�E��� UQ�&G1�.j�26_�-:����Ź0��c��q�������/3%z����G������´ɜ?����Y�ze�h�Imb�
�e�5XV�R��s�S�z��'��rpC�Z����^@W���&�h��3��a\��Qo�O�O�}n����|�����j����`l#��Fg;s�e�o�JDe��(DXE��BԯJ���8�1C�����׾�����>������+��h�ǥi��P�{R�^y啅0�1u�\��� 1 O�KL�Ͷ�)��v�QF�E��2��	a#�ݳ7=�Q�MO�3&��`������N��YB�2�X�Ɇ�\w׏�����p�&U6�bt E�?��?.�jb��Xbm��ĿF�'$�����^���s�={h�~�2̥����ƨh�[�[���L9W���`�L��4�Q|�( ��	}<�~�
���a�s�2���I�Eo�6���7hlv���Է��&��9��t�����O���uY**J2�eN���ۓ^�/H_���gr��slD�Ƽ�g;%0jee)���KC�;���\M!��iQ�F<��,�ɍsL�)��X$h� `�qx�@H��v}qM�#�]?�9�)XCRx�m�JH�`?�ߝa�@�/���xEz�S���@y���9���� X-���z�K^���O�tRa"zV��Dڋ����u�1���Ό���>s��6�K_��t�����yr,��ե�UP�F�P��p\�5�b��DSfu�F����/����
���e�B�-�4�<�����RLS�._�z����'Y'|*m+�jlu={�|#�矦���s3�]7����a�Zy�o�
O)~���	 �ٵ��qՕ�w~���S��t�E�j�H���
��t�+(e�x�i�z^�a��3�� � f�j�pǊ�G`��W_]��
�`m��|J����{)X��1�馛
��}�Cw�v<bn4LFX�O�9�I���?���%q�s#hS`f{� D ��l=���� =P9�ܮ����{�yt ��}(}���ۍ���"U\�z[o�\�B+U���׾"���t����y�V˥�܈���A���H��	Z�6
;��U-T��GU�F#�9$��琨_/�b&�k`�zf8���g|��i-�F��'�m�з���TJh�����ot��x7A�I����rNKKi����[�>��\� �c��ֆ�N&����Go־m�b�#�Sy��J�:�=�;_gO:Vr��t��/J^zA����b�[]=���K3}���� $����Ӌ_��w�[5@H{�;�1I�dȼM&R3�������;L�B���"zd���/6�I����a¨#���w�V������Q��С��y9D=�D���H90����t�;m I����e/+�!₺S���O˥���;jW:���F���oݖ�;wEs9�J��]�����g�9i���q��x��/c��z��������\��j��J`�d�%�ƅVw@����~ְQ��,t��ͲNG;ϣD�{��xZT��bܘ�<Z������77b�"@G�����M����F�q�|��p7������~��<W���=i���]EW<U��� mU������ �?��?+��@L�Ԙ�Ԡ$��T �%8
�dyf ؠ���գ��z��������Q�vm��M��N�Ǔd�ߪr��t����
Ӣ�0�J���������≘��c�w$���~��������=�yew2��:��ӛ�[Â��i3��a7����O~$?ǝ%yLw8 Bno:t7eY�dqk0f�c�`������B/��Xj��b���gdr�䜗�nu�1Z��_f ����l+]������~�3ݝ�h�L��T<�@�b���h���+螥Ǐ�o:��^O�Y�:k�N�
M+�d ޕ�����#�#7|*�������ƹ��O�:�y�i8GC��6�A�^%g�)"�+�>��t�7��X<;����s^I� /�����D�Dc��zt����<��#���O~r���k�{O�O:�7;��Ǐ-�7LG`y��7h�.ߣ��0�$�7�	�����s��a� UX3����ԸP�b��Dy@x�A׻2�=^,��A��[�,�lwW2J�;��z�H}���Dp��P`����cSP����CYYd\����v�m3C�N<{=�JF�/:���M4_O:�]��Cg�9�c��=��!�y����������yMt2���Ez�kϧ#�g"p��^�x����Sk�R����Өt��3aUeJܣ{Я�گ��O�_�ksx󖷼� ����rN}�G�R���g�:��F���H�@`�C�Q�BBQÊ5����L8��Q<�IfЏ8�s���&�Ao�>���6���` ��P(>��3���ท���e��X:�����{�{Kgt�����N���
�u�U&%9�3C�Q�O�!��!ї�ۣ[3�g�|Ƥ=��~q��|�I�j\b����g����1��� ���!?
��V����P��7^s'�7b�H���S������77�9,Xi�;+�u�Y��$N�y]G���:uuDQ���Y:�f�^�ղ4��n����i���k���-@�_���&x�j'�cLpϽ��o,j�c��g?��x~>ӥR�˹�_�
�f�i���4�D۔BL���&�W��6�U`o��`�F�?Z�,�,����������l�UԈ�~3���b����`h��\Oy�Sҫ^��I'�[���N��z���]��a�:"N���]>�Z��,n�K/���ӘOݕ=yw�?�g��#�
�� <J�zz��|��؜@$]��ͤ#�� �A�z�gN����t��$�}:��MR	.����3]'Y3,~2���5ZCD��l�w�D��Ѩ|�����M�fb�����Yo�Uo+uB�Ľu����8s�T��hB��L������g_���\,7�T��1�s� \E��<��5�����t�5�U ����T��?Xm�g׌^��4�=&��:JVR�n|f�cQ\pW��Q�qj	�OHQn�^1�IRv�V��Wr�iD���b�[��s�P�3hQ�Q �'bɯ�ꯦ����(:|����g�z���4�M��bzы�Lg�����-�fs>�����?�'�:��j��W���/� �Q�$�9�>���V#�d'Ϧ��	�,�v\h�?��Û�u�T�
�N��9��֯����1���T�*Rm��Ҁ C�a����H�G������P��������4��/`��be�8���h�jN��ʀ`����tn^Co���^��g��YI�n�v�����l����h��Kq��\�'�nhu�6���/#���3D�����e���7}�zrܢ�>������Q���4�
�muO�7�n�5���kV7�5��wח{l5��x�~Y�zN�ĺsˢ-?��w���\LX6L�-�V��!�b[£R%�9���ܩ��E�Jn�NZZλgcWIFR"{FvY;m���m����lOQQߡ��1�}�p�~����QT���
F�i���ТԶ]��@�o:����o@�o��
�3E�����ck &��1��s��� l�k���y�?�Ò
��ꗴ���R^G)�;�.�i��N^_�y"W�(�����̩0�q�Z��(<Pi�ˢ+�U]1�`8��e�GOu��F�K����@�3:H�� {su��5[�Q���7^̣�I�JG�@FQY@�n$��Id�E�b8���Aa��/�忤�����x���S�{&y�@�p�}?梒�w��]��G�N����R��Z,�s�3%�)Y�ƽQ�xF̬yKl�Ec@l��R��4&N�i��?��(��F ���F��,+&������i�#��?kL[7)�)���[�g�f-���5%	2$��9��"o�����N�� ;�y]3���X�Ъ�Gp�B4�q[��sh��(#&��
 f�*"r�~i43�����8�7�?��R1p3�G�/�/��/n�b���/K�ܝJ5���KH�s���&8a��qݲ����o-�qG�x/j�4��{��__6�?��?�����T��E�UF����Q�i~��I
c����j;�;ɶ�N��7��(�����e��1��y[/*���w��99�w�R6|f�Z	�X�%��������b7gpaLl|S p;_fASE�:f�i��n��_�n�t����%O&&��4d�..h�qhGs��;�����@�Im��;����X0GНi0�`L޽��آH����4 ���z���UND'�[V7o�7~�� s���Q���4bT�_nhQ�S/���@$g=p�qtKs���G�ܕj��J$�)�����.[\<�n��O���7~/����ї]����/���5���R�s��� �e�;�=�)��ozӛ���jbw�"}�Ā4ab*�[G�n-� �Smj$�����)u���	�����/Y�mt����,���=�:���ݭ���CE�a8L���U��������d춵�����L���|�L����7_K��c�׿4�y�A:T�s�@����}I<2S�Χ��f�+Y�e�yY�GЍ%�l���nH��F]�|i,D3ũ��1(�D[�}Ǘ�C_ɜ��1Y
I7Js@ˤ�}�g� ��Cp�XT�1�Y�}1�Y�OՄ*9ƈ�8/�G?�u׵���GԵI�3���CZ�d"���f5}�7�C���y��M�3Ӡ�7�h&1�RH����Z��d������Dʰ"9}������whх�y	Vq<R�D�9+fG��͚��`�5�8�n���΃0MŽ�ą���yl��{�7?H5QxX�G��N.2` �cd,�6>�*���]�c���g��GL$�	��\�>TvI]�bL��ހR~7K���G��_ �LY��~j���=UG�\�1~h�QO�99�������E ��u׶�g����bFOU�=����dT�O�G�����kxV}���KSt�~������y�K�[�$bb�� �R�����ѕ������
*B4���'Ԋg�Lj6f��Z���������轻:�\�2��ۈ����^��i�Ա�y�$ B����}��.}�Z�_�7X1�d�a���9�:s3f���/Y���4c^���q����Ou[;��F�q
���L���z��x�v����M�f��e�WUh�-�����>P���y!�DL�/|�El��8���7��t�'?����L X1zb<30�=:\g��:��,���`�i���iq)�`��=�@z�c&�gH�s�ʢ�f�Ԩ^��S��2���/�7�c
O�l1'(!��[��\� @K�����o3��6ꍚ��µ`�0.�1� �p�_4�>M���`��nP��Ju�lWM�l�����cY�(�l��Ak@��Nj7��L;R��	/��#.97}盇��b8"'L��Ȼ��>�id���ɧ\�Vz��_����� ,� ��9zaT�GT���i�/ǰ�+��`!T��4�G��	hƏ1��p!؅���0��lХ|��0��۱�^�w��~���(a�;��$#�����N!β禠��1�����fq��Pο��o.�9���hX7���-�F�6;�L�\z0��%�N]�_� ��f�z���{q*蘆zrv������C�YZ�1a�VRIo]�L�aEU�V�a"�D}��1M*c���<��s�n����-O��'���p\�HP��{�~ ^��^�xCf`�J��LMu�L�>�m��舭��� ��֔���r"�=��g=�n)Rz��l+�3��O/~�u��dl�I�|�h�
o��TI�k�Kq�:F��G��!�}��^{m��AU�O}j�p]]:}��Ma$�%�C�s^/��'�8@��%�N.���oi��#(�93����ц<��?���{�t�ŗ,�?�V�Šk8q"3	���X;����Iq�1�,nM6��mq�G>�ѓΨ&{�zhL�ed�X�|����W����ͦ��}LZ\>�fڳi�t�T%ܝ<�*#\�3��2�*6�g�[�%��1b�A
&2��&d�ɞNT'�zz<������T"����d��O�C ��������@4VG/S G�!�Vw�aql6�}�dqN��kV��5�� vӆ�T�ek��Z���'y��3�`�V��g\�Ĵ�ey}��3�<���#ŧ�����������I}���-0��V�@y���EE2��&�s���֞����#5���������;�#�ӯ~�u�6�p�����Ύ��^&�jeG����z��/|I�ǗIȎc�"��.8DU����ތ���G>RحF#�TY���/:����4YX��D���v�)-�.����%鬳�(�t[���N+˽<A��Օ�0����үQ��l?���80F2��W�i��f-�" �;��/-���)���ۉ�~�w ��5�(��<�����/��,Y/�!kG]vd�����l ��p�
�	�d�l��j<g-r �=�����:hʹR�C����l/��XI{����v��鑏if�r55;Y:Y��n���k��j��ꪸi�o#j�L����!pT��y��5���y�hxv�XHϸ�2.�	}��a�V�Q�~F�ÆŹq��5�Z�C#�X=��L�֘DUU~�3c�gb�`w�ywȆ���*�� �b#���_�bQn�� ���7t3�~���L8���Q�Ϣ6魎E�n-�����ay.e��a��׿����oڃ<1��مt��y@gw�!���n���+nzD�u�U���PoV���{��aA0A�ie�Q|*�������7��9�\�C"�N7�	�>��O;���w��2F���	b/�k�˭���K��3�p`�Jr���Ƴ���1�[/^f��.9�˔�fb��X��E������' X&AA�eʅ�f�`6[���0K����3�%U�#�����|��Ԟٗ��=P�� -�ߝV{˕zb�Ve<��^!46|�� I�6!0�������4�K�����
!Τ�%�i)CCntd\�_^0p���w�l�������k���qI�CU��7*��X����0꾜:��a�kW�zе���"��q����%ȸ���E����X7���a$ ��濺1���Ci~���*��O���Jlj�˱�i��Rߣ�����Eo@Ft=�FٝhηXbD㿑��N]�y"��^Ի�7���=�O�`gp���@���FBc-���%`	%����u��ArU�l�w�u�T��F:�z;�t�x���D��{����Ꙇ�� �p0�ڙ�\���ff| ��MeW� �������6`�N��7���FĜ���&��aM:��T�5�$�[p ��CUi��O��ԙ��E��������9O8d�\�v!>�3���[&��&�| Ev�<t��%�D��u���ۛ�PT�3 �;��z��q��p4�}�����O��9��Q��=�A9��ü�������
�x�\ԑ]2	g���Dܮ��j$���cܙsQ�|:Z]']7ј�z�0�!"V��l��74�&4#�8�u�� ����%��M窚EI����>��-�G�>��^cl:Yg��]ψ��TUmW{���3��Ŵrt��9X���_��-��/s�V�L$'$���� ����-�;�o6s@���(�<1(E�� �IA)Ƅ<��qyŠ��n�Q�9��G'L�j⍳菂�����swpM�nn��6�T����h�h�����u:��	�P��j\D��������i%���l��#�9��V�$q�lU��A�\1�������4`����i1
�D|��jaEN�4�o4���K��<�Ws1_�����orQ}�C�S�+�3ݫT���<��=�C��=!y��6##�p5�O����I&4�yu���J��ʌuZy]f������R�]��vJ�!g����J#��-���'�U��>T�#TI��FP�n�5͋F_�hߊs=[O�m�;���h��n��\��ϢU���-.$���4�n�.78�fLL;�D��5T�pK�/��u��,B��H���^�5O�cu�-�5n���n�R�c)���?=�nէ���P���;�
�űӛ�;�ft���m��H4�,Vw2��vԅ��Z�Z���)��1��(�,��*{N^��#���6d���F��:��sˈ���gh�����k�K�]rNڳ{��Cbڝ=xg�Ӯ�*�{�y�T�k��g.�������ّ��b���t;�y%�?ٱ��J�FqN���ʃ��{�T6���|�M1MuSh��	��`T�6֘Ҵ���\����J,�W�u}�h��u���&������G���E=\��h)=��'��g��r�;��sF��H���?�n�-R@��xs��19�9#d�Nds}hMvb���vYpl^C� ��wJ�q"��!���4ؔ4~q_|f�\��F�ׄ��t�ENc� . -���2Gn[ �ngQ]ǵP��ր	��@aY�(��&6��uy%��e���=���k�s�{u�(ޞٓV��t<3�]{2;���\���SXtņGE_K~�z0�FW�W��r�(J]p���TM���)��,�.�Ӣ�'��t�@����Iw�N�G}��wu�R���Y@]����ˤ�R���kO���0H� &���Iˋ���=,�<)�ͦ��F:|��#��w��f���VTaT��R�A���ޢ+�(7MdU��i��3T4�L;��]���玢*M 0o�^9,t�$��F��u�ܵx'`��ݤ?S�ZA�y��#�ٺ!a��/�fߨ������G�5�]��/�^�)kp�Vj��_����)�0����J:��FqUC3�j�O�+�t������L�=���cX���5�)��Q�ZR�8���������M�c��c%xu�1�6�Y���{-7��MAx��M��z�3�)n_щ^qJ�(]�Q�'{|/��3���Ȥ�P;�	��J�k�K��>��򦏦K/۟���G���۝Ť����®�<��lK������i�I�PWO�uc���i��Ӫ	�Of(�>O�q�~u���z2p|�ȯޅp����`�F��o����� �!�%�3_>l�	U!���u��X�����6"�h��k����:Y*kfiq)}��_I����ӓ���t��Jǎf��ٕ�-��(����-^��Z}�~ҝ/�O�F�C�_�?�Ҳ�$V�u7ʺ5F;�T����n�:����RS��-��Y�hQ�R���5�s�~~~�e�^;2��ǧ���Z�TϏ�i������t���7қ���~�.�g�yR�������Faヰ	�~$���|V7C�� ��d4ҝ����`@k��D���TtC�'{O�5"��m�2��$ǉ���A��n"��`%�B\;4Y6�|��*�~�<�$̣!��;TlH0������'kl2y�`�:��bجW���g��+�7������}��ON睷7u��|;����'�Z�*׮䫞s$�����9�;��ű��N�w���:j�5rwJ�~S���(ߘ\b|�k�_q�h���q�(Fx�'��,������_��1�zu�s)�=�O�<I�����&=�W��>��%���2�Gg|���Q��x4���N8Z��i��t�<W��  f���������<��w���Qw͹�zy-�g�C��Z�ܒD���Moð���)F� �sN��P�{�X�ي��:eذ�]"Q����Xj�Y9���Ψ$jG�<r�h���8�Z��v/��V�3ж��LN�G��z)j'��>C�=U<��umu�`���D����'8�q<tџ4�Tf|0;!VM��1�Zd�3{��^p��:u��|b�M�RUy��,�u[閿�3-/Qv&�R�S�=Wr#�$��I��Q��Pn����H����.q'T�m;�[�,شE��N�s�r�df7u��j9ݩ`�օ�� f���� ��c����9A��djzr�⼀7��]Y-/Z]=8MT��o�RN=zdt2;˼��b��Iw�u_&7�t�E�|+�ػoWQS�
��-k��N�7Zw�mbE�k�q�k�uf<V7��)��MA��sv�dQ�ڼM��`"�	±	�u����ؚ�q�E����w�-�r����R��f暙)�"��ԙ���"���3,Lx<l�ᜰ��u?tq4�E��rӌ��p;-2���9��4�Lk�C-�պ�wBg��׼�ll]r�����a���	C����bXSg�a�k�� �a�a�oX��Du��wDɡ�`�@%�kZ�����Un�Ʒ�$ٮ�g��m G@���5O��y-�:?(�H�Cz�fk��+�̠1>�f4u��ApZ��>#�����ql$�Q]�mLQ��e4K���l�gQ��-�.*�xg����c���n}���3�����T�k��,#���3��52��}/�ڛ!x���K�����t���ґ��y�P�1�q�[o���w{�b��v� W�nd�Vգ�h\U]��X�!l�EU�j2ϭ�D\n(�\#�ȑ`a[+`����9 W�lh.�h����P{L�8+��p�>�&��I�F?�Ra�|+��g�s�>�wϥ�_��t�p73�R�����JZ��`<[�ёw�0��cp��r3 ���g7��X#1���љQ��wx*lxsn������	�t�2Y�����|ŉT_Q\����Z�U�#G����]�RG��ܮaz�k_�.�p&]��+������r�s#ZM�/�r�4O�S,)��������� �e�i5Ĵ{��	6�	ڨqO���QԮ���4���zO�> K�Q}Q�����OY����wo�(Po�$K�?�b �k�G���f���Ͽ�{_I�����������lvP���ٚ�l�\��4���>����>'}�w����URY���-��J.��z����]�˳ҷ�	�9��a�
�p=.^�q���MAx8h�0��0�:�x1)�Ư��x���6M�+�C�k���D.ӌtu ���E�;�^��̦��ܚ�7�^8�Ծ�$*q2ڗ�7TK�>��|�l������C��h]7L�	]d�&Y����4釶���ʄy�f���}�<��l�uт.�#ޏs��PQIX)C�<���Vu�=�#�9�I/%}���h�,}1�2&6[5���n����O��s��tB>_|zgJƲ�\�����ݕ����Һ���:�J��]y�<��oN���E���$��.}�O2��\�`x�x��޴K�an&�(�`7�N��5"EG��O���/�[��t�f�0���AT"��٠l����h^O|��5�\S�g�'�(͝�&��*<͐T����~�+_O���L�+���);�K�~����6*�\)�R�yTÛ�M&,�g��o������IFK���͌s�xND�y"M/1�Ĭ��ɫb"��PĔ�Y������`�(���d7&׻�K�{%F��K�ϴ�i3���6�^&+�O��̂WZyø'}�K�ʠ|����p.�ʹ�{��t��invO��-���8^��h;����������I�Y���s2���<�a�)�S��-t�Pr�.+!���j�<��^z��W��{Τ�9�2LE+�3������:M7�tS9>:��>c�����/y�����t�UW����-��9d����o/;M�B��}|�����A���[I����Z��Z,9���y"��Nǎ؄��@�DZ�Vs.�0e��P���x�p�er4� A��^�<�����9����Lr��i3�>��O;6��Ģ�3�+ L_@4��i�\� g�,��E�K��G03�}��v��Jȵ�t����B��R�'
Õ��c�(j�Z	�ڿ!`��"ޗ�8�_��{���tÇ>��A��I�wq��OJ��|)������)��:I�d���70���^���� %%�ԛ;M�M	��4�~��+��#8w�7g k0��G�Z�CI$��<-�Q{�h5[�����)�1��,�'�ܓӳ�y]ڳg_��ٱa�N&��x �EN:�T��V�K��V]�j��ԔBd�?���.ߛX<V��X�1od���|�]��d�{h�Ҿ����f�f`����nx46$4�9XmuD�iup3�D�&��n'\��O�\UCXN����t�M�T�V@��  ,N6ve��*ki{uۀ  ���+nz�����Zt�����PE=�6K�����Ozz0��O�ռn��u�Z�MGC��s��u[fó��S�Y�UW�K�Kl-�{�/fD�oc�SQ9V��&�8S\�����7JV�x�3������k�9&����=8l�l����+�O5 ƚ��5��d�A�6>���yIf�ץ����j�h;1L@����`�щTL%3�ᛑ-��#�9���`>N\��h� �3�peۃt�H��bR^L��2��8��9�x$�#L�1�-7�J�<`�n����n�r�	
�7bB%��E)�%�j�ZQL��+{�0����^��Έ�6a���(�\�����8ǔ���0������?��-",�Ρ8m��lR�W=��'���[�HEs��H�����3N��B'��%��WRZ.��о�v�=#8X�a/-����[�y���+éj'��-�K���������x�;J?�[���CC�M�o�q�4jL@L"�9�U�P�tp~3F`�VQ8�͕�v��d���i �����~#?��t�W���~=���3�;Zyo��I�P��s��-�Z!��>�/y�K�w��Ǽ�u�+���b'�X��0�z�	�$�LN�����GfJ�~��-<����S+l���TJ�4LH
>�A8�t���I�	u�y�K�9D{栬PF㦿�0M�\��y^�E����cX��0�EC4��ҏ��wu�y�GI��晽v�H�k�Ɏ$��௚�r_���V�r$]x����F�T����.ܥ��<&u����/�{������ )�fc�!K;}�ӟ.����P3��1�>�&��� 5�;*��1:ڊ"��g�������1c���}n2��N���h0��/�,t�W����)`�t*`�e��{'+��Э��2QM�����:)asF�=�O}�:Jv�v�Xz��H���I���4�����ݝ���/�Gjj�	��!J�V���|����{؉T3>��殺���et��Ǩ�nX�fF���h�Z 0aĬ�]�ۚW���7K�RSVE7W��Ut�C��)1'�a��sG76��Dl��Z	�5�܉��s��RF�f�iv�\z�/�<����N��^1|�;s��qX�\j7����uG+�_���n�ES�B5�A�1}�я~��R� ��RmK�q��� ��
��>�s�^�(fx���3
 �G�h���X%qzK����R��L������!|��a1 vI� 8�BG;���� ��yk��s�k�oD������_ˠ����[�^L�������<@�i+���{�&��K���RvTJ��Gm ����H �0�y� �9����3�h,66]Æc����s�噙��!��t�YG�M��:\�M~���]�Q"�𞱁]z,��F!H�w��r�2��N����]��^<v��/9��~B�������L:v,K2�nI�ngf��R��y��ݔ&�rm��7 Q�#ρ�FX�)��4�0�h3�����
=�/��➼4�2���ê�X��;τ�VAv��^p�y�#��~XtK�nR<�)�5�#D�B=1��,s>����ꜛE�e���zX)_��W���J�]�1@#����X1��=������\zFz�k^�f��<p�8_��I�L�s��@nϰ���EO��&[cc>���U%�x3���0K�u?�m���h�tB�l��>�����@+; s�z��u#d�3���"F®)��ҪM�T��y�7��Bj5��K��0�/9��I��,5馛>�>�gQ��ЏN�3����?���l�uE!b��}G��׿��E%A?��.�U</�y�w��]�>%%<�x�3 �/�P�Mi���Ҷ��8��q�]C(��
Z��q�y�s�����bqgh��}��W�� ��Ibuc��T��xH�-����B���qC{�k_[vA���t��t�;���"��qq���2�.��#�/��>������;����oo-�r���L�1�e���"��DܿO��Qׇ���ԍ�X��X����I�J�,�t=&;�`�Sl�ޢ��{B�C2�'��em1��x����~�1�&M���;�K�X�a��fܞ��z��L��+����=���_~�3����ҡ�{�7��t��{K��fs6���R�3>-����y0ȿ�e/+��.��oxCynt�|nE��!�XHb�b1(��(�sn�EyN�Gm�=�G������ڈ���UG4Z�ҵ�[%x����$���ۀ�$oc-��;��+�1������"�y�~����������芟��g��e�q������¤�sh����ӝ?�7}�O�:��U�K�>��H�b�+j�F����Uʲ�Fy�7i�Ֆ�"��XMs�[��m*)���&���b�N���&�Ci�~ΓY�^G�k�s�qm� '�I£
�{9���K��;2��
�3�%�Xa���`�,q}��XŢ=Eo	����õ$@T�"�a�;��owf�sdm��U�������t�������aw�u�T�f��3c�W�,�	(�̪��G�e��������˛���"��;�,+��������x	YS��O�~�����S��k�2H4�L���8����'=��PG�G�V���ʺ]6]���k�ݍ��S��dwٲ�_d
ՀV:a:#�C��ab���\^ӿ�ɕ돆ie9�C?�/��<IF��[�H�_p^>���� =��\�u�-���+�? � �Rg�?���.̦?�fA�U��L��۽׺��k1_�/�L#�� ���h��4�kØ�7���r�fk~Ƞ�E�,��^�}��Q�,[Vա�� A��D�M�!l��WW��J�b���]E���݇Ұ?���ޔe�|��������\e������7� �w�H�آ�J@����'��5�)nk "�D��^�)�|3zOhP��^��	)1���UQJ�4Wv���R�hT��/4\cavRw�f-��."ѰJv삈I5h�υb�c_�җ�����I7�pC�\X0j
\G���?���"]�y�oa~&���H�>��tɥ���fz��}�J���+m�����yo�F�>�g�����:ӭn� .8�n@�ewd0��E&b��9�ew;´�[��
���Pώ�z�-��c�y�v�q|�<,�A��xǄT�SC��W~�p���O�_r@iD_�6Qݻ�s��\u��<R�k�Է'23l�Rg��.zę閯ݟ�C��WJD*�#7e�Z�̂���~��9�x�$���7��<�9�?���T�A�~���wxWi�:q7>]cـb��8~q����X�X���W̭���l�s;��h��y��r*f�|��z����;o�ܰ��sx�)ylԁY"����������$5y5l�I��|�3�)��23Fm	LS��ưL�QZI������_|Af�g�W�+CIU�QXq����vU�S@$~�ӞA&<���T��fM���YwK�Qb�m̱���T�a���*�#�ى��F�I ]�̀  �� @��)1���[�.�c��!��ڊ��kK�aT�`��QEp?H�lJ��j����!�W���if���ϥW����;ߺ?9�/u纽ci�ފU.-/�
+V9\��+V;���'�X՗����o�v�P�oHƀ��싸�}x=n4���x*�4�����}�mu�E�b�*�&/v��@͙�+
Ɇe���Z����g1�E�gXA�F��D�<�'�����u�G}w���)�Y<������t�#���_qQ&�t�b�U���**��J/�~�f��6��D�u�0�L�M�)����n\��N�im��4����U�O��{���(��J��!q|��z�H}.�D�DI�s�o�g���Q��X-id��2�<n�[��/�a�f�XmF�6F���C� ) 0��	k*��}�������e�|.�������͡�OOzʣҿ������Ng�ufa�Ԥ�u�a�_ȼ��p�IG�z^?~�����/�R�PF5>plԑ��Dn��TS���Iċ��Qu�����d�����}#3��p0� ��A����shb�b�1�4�ޱS�!�L�Cǘ�'2X�75�:6un����uT�E��;*�|~�0]}���}�.���X��Υ���i��?-�3#u����q���6N�=c��:˵�.�N����f�Fu��'{�h�ޮ:��D�`��+�v����國sW�<@�8�0b�)`k�M��vp���ͺ@#ܭ`aVW�	���_e���fL�!�s��@o[�_T����iFs��������˳s�t�Ż�Y�^�n���L�qSg&ϙ6*�n��y-���R��0�=��O��C�����Pb��sLc���8�Ք�ԙ�;��6��&��W���y�Z��E�q@����m���F�v���0��i/z����+�t���ID7�>Fk����/f�ѱ��7����Y��q7�9\��E� ��� δ���}���T�$:gG�����A������-}�;�����M3s��޻���eί���/����ԊZ��@�iQ���+����K{�n4.x\`������������4p����:�Ό��.m���ν�U_��A2�Q��	��L�f#�dmH� ����Ju����m.c��8,�kFC]TM߀6b���y��3��D��k^߼��t�_|=�gKY�Ngwcj8��Rf/--Ri��:YR����fSM�S�+=����ځ8��~d�yғ�Tp�M�d`�Ȍ���Ȳ������r�ʪR��$��Ҋ�B 	#$�	!�1k;lf�D���3቙��n�{"�1�&�=xŋڣ��2b�X�&�RH�U�de���߹����n��r�L$���Ro��9��?��1�DԲ�1A��zL��Jrw-�asc��T��v4�[et��)1,�D`�+�ޢ�۽`�{��Ŏ�������Wy����L@���F�dI(�tg��}��Q�#����
�ӟ�L{��L��¿�@�8��}���h����/3w�Y;rx�*���E�;��7��Zb�]���s��(5����yc�6!��� ��Vmh���ă�V�B�K o.���}��7v]S�y,iF��3G�$(.��LR��浤DU�`�(E*�6��������w��W���wJ����pkAj\�}���K����LP���-��_ ����	ϡ���ȋI��趕3Yx@pUL�����?�~#��/�R��ؐ��y�5�p#E���g�
0��_G�)���ø"���F�cUdֻ&�u�N��N�2<�Z��؅0������;Pc��i�3qxϮ)[�De�(�D&U��N�k!�q=�0�J��@�
��#��2����[>��:'¦�C�?��V �r��ӧ���O�f�`�Y�\	s\����K��f�5�d�^?�@=HϹ�+��_�^��u�RE��T��4��ȧ�	ӭy�C��km(\
D=��m��@�����,��Ԥ����"� #n?��|�"���"�6�÷��.���3sԢ�N;�jVo��|���frpWm���|�*�}aN�D{K7���+�^��\W�\��j#a�������g��0b66��J��ؾ�D<�P������g��+:��W�͠7���8���ګ#"��$fg���ِ�'�z)B��'í�!�K���L�Ag��@���X�M^I/X��r7RzLO���&� �$@��85�OڲU�jV_���#ǭ:1c�V�z��v��@�2�IA��D��p�C�\�QQ���8J<��_K��:��ꈥ����leD�����d�S��S��B��Q�{��ET/���6�ݻ0-#� ��}bڎ?a����rXS��%o�	��'S(�j��i�c���*:��a�b~��T?ZK��BlvHҤ��qc�C��y\�{�H��s �T���O�6�|<W=��
�ЩY60�sQ��N��k,��(ّ�XE~u�
t�F3�`���X�Y]�^�Ʌ���|gO�-'v"j���:�!��e/pK�u�7K�L��'���UJa'���!ڝ��}�f6��Õ�9;���?��#�:\m>E �6��>J_��+�����J��L�Z3^�/0՟���|//-��x� ��Bja�.�>�l�Y8%��|���eo?�n��%v���5�#z� �Y�I�)
@'P� v#��<Y�|`�����/��{�Tr�
9 U(2�-!0|�Y
���RܗvQU��<P�XC����W֨v�$�^���I{:�r���ZqY1B"Z��>�������_�'q��\�zΐ��@�K���޲\B޻ m��@����]��a�hu欓�;x�����_{o��ɤƦ0�[Mc}�,:h5$jM$����������a����К�R	m ���rΫ�._�����z��h��>�e܉�O[��`�j�6o�loy�+�U��>��k3��T�@��Y��rS~r�z+%�2f��e��sA���u��l��7�
����=@����x�8"��:Nc��2/D�����*�ʟ�&F(��,�m�\o�s�O �Nf��Z�bZN�t�dgR�W����A��%��x�(�׏ϸ��`�Y����Oy�=�'Æ7|��1	b�FY�];��J�c�d�S[�f3�n���[��軒Յ.{#�!Gq1�!|���a!?^�"����(�96h<�~	x�3�j5��rA���m�<k5�X�����42����~K�[l߾zn �t��@_c�&�����20{젚��^T��� �0	���SQ	�U=t�✹&@�Ď�^AJ�i]�������~
�N'�\��70�-��kWzX�ۄd`P#�������yp�� RM����T%x���lI�A��B�n������l�[n�:습���v���WZ��l�&vx5���݇��Q�<?��w��Q4�h��9y��=s�{�]��=AF%��ǺQJ��0�[aݶ�6Q��q�ngE�x����W��]q�Kl�maΕ�L� uv[�Z.j>�G��(�P̛����9W�DEo�(F[ ���q�W�e,S�>����6Y�`/�&]7l���p����jt����A��~/ZD�����-��	<|��>�Ĉa�P�E�����}Z���[��'�x���w�զ'7[�r4�6�<l9��WJE� M4���\�0���?�/��V<�sL�gi�Ӧx*�ޜ�?�Mb9 X��d{3"�z��A��Bs{�d�)��v5��i�����J��r����ޯ��/�gs���_�2H��1�p30s��Mo��n����&)�3!^U�DEb"���H/=��5ߕU���1�:����=��/�^�#!�ƒ�-2�Ҟx���GK��r>�8A�*�����Jr����b`� �{
�}���&s<�[�m[w�S=i��������ο��p�J�̇�N���CE.�G�y#���'�7��P1<�/B����s��h��o�ɴ�EYW�zf�(�X ���"������e2es-�]T��̘� `��>��v`���n='���/b��S]R6�����^۽߭�Z�&5�"D闯�&WL�_ᑷ5q�2���^Hܸ���=�y�s7�k�.U�>މ7��jJ$�7�sG~��8�;�{=�����Hw�c*��E]�o�~ǿ�ı�yX2e�����_&I5`������ӵ~ވ�j��J���@9��I��z�i�������$�C1��O�q��j�<W/	�or�7�&��U��B/���@�Y�7h�o��"�� .h�X�_t_������'҂�����W�)�iX��\fv�ZSv]�*Q�011�3X��^hԛ��Oe* �YX��ʞ�d��_�
@��4wG1"а�?����������=��Q9Y�U1��I~2�z�Bq-���������/��}8퉙8�ʕ�.��۹k{xo��t��V�~}9��"�<�]�[�=��O~qkg����{ ��{Bxg-t/�d��-N�a�i?a�!Ë�:��j)��_ۻ�s�ħ�/�G?���`T�t���W1^��g染�,λ#zfE��v����E���Q7�'a��}�;��Fy��/8���^��:1��j�
�����[�;�EXj�+���Qs�8��ڄ<���or�I����,pdE.�����Z�IEU������{&�ũ=}�i;}�6{�O���\p���(���u%�ig�o���2�[��" V[��P��s�꓀ƃ��"�i<}ٖa��Un�=��Kaq��f��C�ߨ��B��p����"��9�9�^>�gy��1}���W�U{�$��o vo��QHs�?{?��}nkKX�[1,���6��6��j?��[��~hG�խ�:fI�a�f%��$�eU����W��=ޟ7L�YOZ�\�߰�S��r�=jw�R�k��5�c�up�����;��sv�%[�y/8;L��(&MLe��-���p�J��(2���U\�9��yqT���X/���_��׵�3�F3��},r��V5>BI�F��g
�;/m	��o��R'���6z�H/�K��P ��`��I��W�����"�΢$�LR��jiZ�� '� 5�L���y��߿~������y{Ίf�y�! �i� ���)�Zq�x�f�r�.5Ǉm��1�QHcA��rF2��-�P�IQ��5���S�m�z?Q�����v�i��~��sΌ9�X�[���U�����Y;v4tvi,	�X����٢�������@�"Ǩ1й�ĮS�D�g���^>ۛ^���{q3� z^-N�Q.I�|tm���;���{�aݛ�DG������˟�!xc�f��]	g��� u�R�)SB��n\/�2��Пٖ ƍ�V�{ٕvڶ���ө9J�g#�q�,J��d�5���Z\�K6���AK�?�v���%#�hʸc��R��*Z�}���P���z}�?����そ-�,J��a�}�DԋA�*ۉO�7��7�f�UȎ��r|M��e'�fƾ=ŅU����1g4+��8*n
zv��w��O��^* q��+��7ho����?k]S����(��{5Ű>�;Iҵ�;IR#�;^}��QR��&�$!���VQa~�VL_����[�,��=��>�����֌I�[��"�N��ju�QNia!l�]���������_��r�Z���.ُt0��r�=��T<]!��NfolO$~�{����b'�J��|������|��B\U�J$C9f��sv`5��Rn�"�S���}<�P�,+��Pa��E����K_����}���A��V䊼�<g\��.W�T_4��,j�{�N.WV*ZI�>
|�a�f�5���>A")r�(ɍ�L�GD��z8��TT�����&�K��J���I4(�����s?r��ү� Ҫ���)t�k���A��aR]�y?Ӫ�����X���i�gp��⮏؇>�ak��Z�bڦ�7�UW���\p�5[��)�5�>�w�D�a�����U��8�Y1LE��4�+�%G +�b�_2y��{Y��QT}�W/����@�pjo���!����ჶ0Oٓ�0qjv����z��l��C��o^I �e�n��D��$�E}��d���s���< �L��b�J�_��m����< �"� P ��r����W���=�^ �$D� ��|~��⺤?����??r�@�������ƈ���8s�~ ��e�+�\� K}�Ky����RO �ܟc g�!<�M�~��D���򒍣����D���&lQ�09U�Ns��	\/Z̪5IY�mZ����=}��0U*fn<ƭ�s�Ԧ�S3n�8R���o� �MP�N��J(]%j��	N8)����pd]O��"�V%d/�	KnT��0�8e���l� Z�<���x�x p#*�B�#�|)}�>H�H�I�3�Q(Iw�1 �<����v�B�bY� �!���$} �'�61�C�u�^K� �~��u���.5цqEu�(Ւ6C�K^���o�̓��92'8_9 ������w�7%�`���"�2/�@"���k"��]f��}+�������L0�h#��h#���+���6����?ǒ��{r,� �	k�{2wi3k��Tƞ́$2 k�q�����_�r{
������w|j4~����uJ��a�F7ϰ�5լ�ZxtSd��j��kA
	��MQ�#KE���'�c"��j�y5�E����E~���}}���>� �+U$�}�+l���)V��><#ի��t��X�u;��p,;==K�3Q�<I�(&��_n�^zi��|k��`�3AI/�����n׿�;"xS��s�+��"r=>�`�Dz@��E/z�IA�J�mǎ�0��m��CN�(�M�O����7��3�ѵ~*˥��W��O�FLyOx=����|_�qC�TE@/�CWCE���g
�3��c����U�u�ߜ�Q�X�w1��1?�r`�q?�x����[����7P����CF=y+(_,m%/�R�z��P�[ 5�q]@S��5�Us���b� �!�2����e�P��,�	��)R�E����l�36���X�h"�&lێ-��+/����\km�=�0��Jo̕��3	��gI��T�����͑�����G�#�LT���K6=*� }�I{���:TL��Vj3~�G��E��讽N�RIڝ�M���'����n��^xQ �kbZ80�k�d�<&���&zB�DDB&c��B�g�g#�������}Q�p�7F �a ��\�EḰ�� <Q��^����D%�Ī��Q%��������3����
���Im��~�?���N�YXԅ�[�i�86J�Q<�$=x��]!�S�aj&�=�L���	�c�Ј�,0/��V��H t�|f����8�9(�8�y�F�25�#��1��X��E*#�a��\-t����VF/Iq�Q���y�C<�r�;�t��}���Q��aé�r���2��܉#�%aOڵ];�����F��/��Z���0��Mx�V�Z�6=#�2�[����I��V�4&��+^�
���ۣ�8�ӗ���1/0e��z��C������|��:,���4���x���Y�<�����v��),a��M�,�Ns�n>�l^t��t��ag:�W�
΀�!�p`�Ʌ�]���j�}�����ʎ��"c����Q��w�i?��?o�''+��u��H�-��h�����ݴ�w�<,���/>m�f��E�jŹ�>�F=p�)���֫5�u�^U�d4!5h����NznΨ�5�����,nE���s�3��� ̢�w�ׇ"�|q&޸��<wDI�f��X�,�é>`�����.d^�^|Fg�x����u��F_�I��SqJ�bh �J��A�h?��E����0�6m� �\�)��?sԵٙ �NV���F�c�[&�3�Zu"H*iۦj����M+U��Z��e`�ݾ;$�P�UkC���������+_���9�o|�#C���I�>��&ȳG�T��넥�{�,��!�0�G ��Z)�px�k�	��(6��M�͛���l�� ؝��yf���	�>ɧ�I�?X{:���.�"���R u�kq>0"����ܱv1_tO�$��7t9G�Өpן��sׄ���l��M��Hy�p�q�y�r"�[=��N��0#����H-�QRzMMl�V�<�Oj�0���a@�O�(�PŰk��7@���b��es�).�k�P9��ec���9ǵ8���5�
��\����yϢ��zp���,\��p�p�������%��}�o='����0�5N~��S�	j4�1Z7m���
���4�ԷT����߶˞s��>繡�%�Q�+�$�����_�U�!�C����s�p�s��%%�o��Jq<c+@FR�馛�3a��5�^�%FI�<�c޾�/������/�g(}�����%��������&���9�X�ͯ?d���ý^�`Lnu��G�k��6.�,nC��{<�������|�#��?��?�7����Ap�StA�`�]����:e��_~�����oٿ��_�߷r���|4ט(���4L� @�B,�|�m�5�G��a<�4P7�:r	[�3�rh�J��\@J�x� ��yϕ�����g�J���E`�$��F��@��a� �Ap�0��o�}��ĸs���}U�$�F	�̱0J 8�7��b��pq\��dh�I�+ΐ�2��8�L*>֟�����$L"�N�n�#�Gn�F����������{���j�˿��&'�m���"��������$�Vyn��u��W��mx����'���}�8Tm�b�Ĥ��c�d^������u��'H�K�bs��{����VXop�k�����Q��������"b�1�i�2�h��XJ�"]��3vFO��f��Q���ɋ�C�̄G��7��w<����"��t�ϖ��M�y�t���#v�'ﵟ|�+���P9n*����fä�M�Vޏ뽎S�n-4�>7,���=�z�azY��E ^Kf8ԟ$�le�l�SD<t��@%zz�"�1�Ƙ,��A�����\��z衞�!b��ay!��l	�7��g�T 9��& * G���Gnm*���K��fA������c��J�����s���稛�Ƶ��n+z�;ٸ;ڱO}�s�������4+'�Y���l�1�5b����?��`l��/��^��WG	��t�a�P�s�=��s57 l �b~@|���֐rxh��yހ�7�7U��P����a�	H�ؑy2LT'�.�{�!��3���#��YF&;��/t�I̎�N�D�a` �{����4zd:����_��x.��E��̊�;>�x�ĂQ(v�DÞzr�]tɥF��VNx2���Rf�[f�r��񐨥�#ø�a���)�P�/��$2�3�@~���R�9 ��� Wɜ�h"j	���3��׼xj�h5�2h�!	�4�>_5s�{���7�q�=��I�r���K�"-|��w|���*�#��!{�|���q��~��:>P�$�>E2�J�)1?6����$fJK����
���u�)�I�կ��??/�O�������8Ό��-�_lzR�ȷXz[ ��Fg�f���o0~y5�X�3|V�E�2w��
a�k�	'�r�M��	�X�t+t�"�GG�k�B)�(�Cް^'H(����u������-�qD8�l�z
0���s�uH���=�)����6�NY)�����n{.:7�T��V�\�ʢ��tn.�D=��* ����`H��wYS;�G��-F���������~�^�Q�;�"�2X�T= �`?�R%� MZ�s�������@T�u����	�5�l�"����B  u��@�W��j-x ѫ���ŤDޯU�О��5�s뙣0��N��ȅ0|[� �i&�����OX'��|c. ��L[XC�6y��ܐ��m���*�:yI<I�P�T$�1��JqTr��v#y��j����ل����J���	C�i���k��хl��YR��N�T4��Kc�2h�J8!������G���:�� j�c��B k�ypF�R+�F��sv؏���p�r����=�U�������D7j{1�b�������yė@g�ܚ���3+�L�mY)yN��?f��kMî9N
�������N�F�v�bëE`�����^y�=���F�4;|�`�/��.���S���0��,��#�/���XI8Tc�(�$oFa��d�+[æ�C}�6�  ��IDAT�{�jS�����ݼ_N8 �8t9���[e�G2����h�XVj-h݂�ᢆn��[o��	_��1�NZ�F,�.�M�Atmj�do����=n�+_p�M̴�Qϸ�Nhnti�p�#R��'��9*m�E�ٝ%���!�sJ�@U . �$V���=j\�3��Î�z����\�z�0�|Q
7�0����n�C"��+i�!\J�����_�cs�;v��^h_r�=��&gg�n"��U��\�U?��i���} �ԋ0(��N~�#�$8�G��! �^]���$n��:FҔ�^��Ͷ·N��ˣ%�m�5�Һ��G�����@ ��7s����� P@����G��N�k�1�<<)=4�HK��\���E�{l.j��]��l�.6�#v����n��a�L����yu��&�KDU�5�"?Y�ּ�B",˫d��s5 ���Z�"�֥���~����b؞
��u�Q��b��:ܵ%|�����a=LN����a������mێ�;�[ϳ�~�` ް��Sf�w�.y��֩�\�ۆХÄ��o��0���>�v�0e��B>�M82�z�(5�����z�a����n�[.-.�xB��&β�A]�:#�_�ThpQ����������K��p��{�[�b����i��{���g��6�t;�|?���|�R;�[��������a��)|��N�D��FgI#l�$@+���Pz?/�+��(�k\��B���*ǩ��Ѩ�4��1~W���{H��c~��+w��p���@�dڴ90@Uk.�b����}���Y����?�J�6���ێ�B��wZRg���|��	k��s< X��{���{��8E4�ە@@�A.i�� o�	�e��Ƒ��K�Nw��5J�v*=G\i���v��¾3ޥH@Z�pQ��nG�uL�k����aN�~Ǻ�կ~5�������Q�|�3���ǃpֿn����_�;v䐕*d|j9|�m9�:s����Ls�\��H(��,�Ч��n\㢉(5�al���Y>�D���E��ն� <
�W�E�jQ�����b.~�/�� U��%e[�_�|�c������8d��MdJ�b7��j��Tmr*��0g۪��/V�2^r3U�� F\$����ߏyq��-�H�X�!�&x�Q_�ˋiz�K�R22ڥ,o���I��n�V��XQy#�h"��:�E����x7o$�3.':ݢ1�Dˑ�G�O�/L�b���3(ɱ�J}PKc�σ�f�-V�$a"a<(��<��Ӯ�a���9g\BU����ë �,�q��ǥ/�q� %#�Oj����J��aTԉS?�>+1>���j�.v9���j��6�g'�B� NNLe��e�I\A��R5��n�gm����|�N�~��̐U�eR^bY�BI�a���d��F+\�X����C���M .�_p��3C�Ǎ���KF���q������{��R��5�Nڕ�#�����p�sϏb�	�%=O��_��1*@C9\��A�NGu�)K��irD̡�G�Agg$���g�:I���V^?]�K�-P�_��j�H�X��Z����J �ސF���ؤ�ܘ�Ae�řӉj�h��o~�+��-�������)�J�s�Ji�Jf�x����(z���&�Fcr`���F e�%Ҙ����T��~������%i7�7�W��>�ASSS�Q#X�w±pɄ����������~�5a�̎���XT��{W@��9C� �|0Hђ��y��-�(�BZ�M<n<55w"�.����H�� ��=ј�n��%�����̎�O1���:��D�d�#a@��1�	���5n+<��ﾻ��ɷ�{pm�����p�u�f�b��J9��ɔ�����M��C�	�K��W�f%��C"���;��+TG��{*r�Ec�8�wW�T[ƵkԹ�8�����h�x=A�_"�&��e��d�sRH�KO�6��8�G�ݳ1�?W+p��#>}�v�/��?�Z�;�
��l�MK���=�	n��{���Ђ?��?s�p�hH�G�-; �8��+�/8�ڒ�?
��:St�sA"������6���^�F�N��ֆ�$�s��2cO�����^���Fu�SO����>���a���� H �`��JN�Ί~"<��?��?�����ꝏ[�|#dD<�8!];&�ڊUx5�r+�؇��]ĕ� �͘O�r-���������~4�C1N~`t���a���n�=[���V �e�6{�Ͻ�~��o��Z �:�Y�&�a}&��%������E����N�5��;�w3�E-b XA�ɢF�@����%&��j'�va��سgO�d�/� |P�����R���3DFGp��Db�i��^-�	�I�XF��$��:���c�Չ^M7���h,�T�'�T�$r�:y�]��^٬C���[b;%NhW�@��A�c٦&7��][�J;2�ɠ�8�<� .��Vb��aI)��6h�����T�42@m۾c��s޶�VH_9���w����o�s�6Mo�)/QS�N�*62N˾��pq� . ���uWK�T�J�$��WG��^�
��ʵ�����w��3�( ��b�b�Pn�bދ��r"�25��dL�sքƱ���_���z��#Gˀ�FB����B
��X�6�T.��蠀����t�ܓ�Jގ�T��+]��q醉�==k؁��ؾ�����fw���љЯ���m�����a�V�Ֆ���O��A�σ��4�ymCkY�q�&����ڷ��d`��
�q]S�sj����/ ��>S� ��T�p�bʊ�%U�����6@ޣ�p/WO��&Q ��6�?���PR�3,�'V	K����Vo.D�����"G���N�)3(
�``v+v!�F�w�*�Ă��ك���׼�78��2@�Oj�z>�ם��Ժ�m�|�}꣟��O�#?x�����ض�;�`i���M�;��,����l���$��X�� �Z���\îҲ�����7��v�������v���ע��4�b�����Ի�*��u�]9R���J��J����� ļ�������B�;`^!��Yد����Ғ �@�)2��-���H�tsp��P\�"�a��v���9%�� H^9�F��
�O�B ���Q^ �{����6��'�x��򃟴׽�v��=-�GIE8�wx���E� ޠ���D�i*�&ʹ���0>��O��s69qF��b�2x��,�� �:�0惫�//@���4�0�!�D;>�I*	�����&�
?1�ΐ�׆��5�R).��h<�Ԋ�^�8.��U;�>3�Ocu �Vɪ���3�C���2(��b�xQl+����������@. UjA�, JVI��g�*z@���R���V���{roVl�����ٌ	���;Q��A���r���ј��Z��o��������c�nٹ�LS�=�q��R|��ԕ+�{H�VjD�2�B��T`�7��W^	~$|.j>s=��Sp�H��ʹ�
�����.��}n�4��>.u@�\NN,�̦�x��b'f���є�V:9�= [t�@� aY�"qB�t\�xK�C�1��AɿP)� �W�|�'�*�z���|Ĭ6�Yi؅�m;N�l�S��ޯ���)��ōN;����ڠ]DE\cYǋM@2 �T%��-v����_�o�*�^�lW��B��^�1[=&/̏-���*F�J���>�X�J �+^�n�a�|ДWcB*X!X�}r��֞NZ�4�#r�t�U�([ϐ7�@�H�G�x7�������XY6�ex|>
��j������O4��w��t������ُ��z��2ʦ���9�T�F�{��h�c��Sk�:t�<�6��r�>����҉k��X*}^4Lx������#�8����+�Sc���}���?�$-?��w\π?6sIMJE꟭o��->E���[|��L_�NJsHY�._��V{�<�k�0��}r%1!�̫V����*�ʡ 	Q^GR���)l]��x`Z��گs��y�c��� ���o���ਕ���ݑ��LD״ޜL��R�+��杘6�&�<��Q�����1�L ��>�s��Џ�;>Y�`�Rߓ���G9����,��8�-�[@��V� ��xw�!4�p�/;a�N���[�KΰK/=�&�Kv���3S5�cXr߻�%����DrX��F�o-7I��W@L�ߚl���&���姩��r��Z#_j��=�H|���r q���ʷ[�ڐ6I?*䟵 �K>Z��_R�(O�����;��RV�%SH�.}cqS���}qU��6IH̊6X�]I�z>>$]�D�/%5��R����7�{����͛lbj2���\w����
{������3b�#\:kթ�����w�����*Z�&T����
q?��m_iE�C�'�(MWǍ�>�����/山��a	b��<�����	9�m��l��Y|�v��������9�7��2CC�'�.�W[.YV[��J��>���X���.U����xx�b��B�X!��6Gq�R'	�]+$T\�mD ��8�︎rp=y���(N�K;j���|�ө��F_�Sz?-lq��bf.�y�bD�U�C��,����$�{��Ӹ*����K�.���a��E��j�/4cy���b��n�풋ϳ�]fss-k�� Y�H���kw���h�h�9��43��+!yRx�P��J��an�9�F��	�;&{�Cn�}����K����&�v2-�QC�������M��i�Z���>:g[gϲ��<1��sP�#N�W� �}�-V��L�,�Sq�J$.S��D@ ��X�ճD��-p����%���(#վw�����H�Tj3��i��y�R�S-7�kN���j���ࢴ8���(Jn}�(4����^��D�}���o�z�r���m0^#�Z�**È��#���FO�jeҞ�7g_{��<�0�l��B7[703��1��Z����3�Tb<����o��Wh� �dFp�˹�l[?�[A��Q;��Z���RWxqP �wT$5�|�.ngs'�W��v�:h� Tu���g�D�F�'7e�"ba�NLa�Df8/���*	)����������1Y<�Q
Pe'�q��	I|g!(���ŕK� (��W�G "}1�䪦"qO�*ݭ6��A{U ק����p=�)�c�VMqഏkpm~�]��~�-\[ܳ'�M`��Xc+���zR�����1��6L���b(�����p�R6�N��@Kܼ�U̢�^�g�ev�;z���߹�����4�Sj�I;|���}���u7��]gY�4��b<Ƣ�/�8�� ��y߼$뙸�H:����\n�9�xUߊ��'��������M���vs�Њ"?f����>wb��'�:Ĩ01�h���	 ^�n���s������	[?��~� 	���cq�X &�^��^�X�8� *�-w 
�)~�J~����$�^zit�Q�@��K!^/������x~���8�w��{"�����M���{|�rJ۩���'ek�$��]ʅ�爣�t�RPEW�� �#��O��v��2(������n�#��$ƕ��MQ�p1�2���H��u�;!���>JGK�i�*�r�+��N�6	t"��"�h3�*T�gGpנ���2^�햔óճ���I�6�FN��X��^I�U��'m ���{yھ��w�G�.xS�Y�ͨ#�:�#q�^�(R�.?�8�w�%^�9�	\�{�����5��sZn��%�T������u\6�S�5�-kwI��-��0��NసVu*��rFT�]�I�"���ʑJ%j���ű�	�Q��N
P�  ����>�� G\v�����ߜOi�����+��"�/`��v���  ~�>�`�� m!3ɺ �.� Ĺ��`M`��T��K{9�� � �r_Tuc�����f��崝1�ܛό# ��*}.?S� ���r-��f��f$� �6����@9�񑏻���w υsy�<��&b�1�;�:���z�$��� @�b�3�����G����9�TX.%�N��2F-�AR�&Y��tлD�J�3ʯz��焇q�ˡnw��	Ot:�ҞRO��*�x�b����E�U{u�#Y�ДA�u�]�n#N���;t`�@����dح��a�΍p�ˢ�?�<�_�D���Ćdܒ�	�L�Z�3�� �D�X�$,\@���x�c��NΉ�R% . ��� h�� `D;��-�K,.�������m��s.`�m�x��q-H�5zv�E�JWʸ�+���u�I;��6p]ڦ�d�4 j���6 `l!�9%cýd�U\3@�̹\������fD{�� ��OWc���<S�XQ(�TO�������`֓�;b�S5k�p�u�<S��;�0*ktӆ�_��g�c�\}����9���uV�R��D_;�	R�TORE%�Ai��ԁ^R�h�@��ƌ�n�B�wB�b*���muc"5���kAIg'qKzE�(�1�<�(~ �u�� H`��`��y\������9'��J%�햛�cS��z��&j%k5J��ɖ���;��G�Y+��="�Mn���W@�� ��{,�0u�҆�Dn?�;:�K�'�����쾺3�	��BC!�ø3�(s@���9�c/�<+�hh�D%��$��Y�� ����/s�Ϝ�=�N� J��xp> H[�tʊ����q�@��sƐ�܇y�J�|T2���U���O�c�#��VF;qb|��*1���޵�����C� 6>�'����G�.���).	s�����ǣv���so�I{�-W��dhC�n��R�[lrb�-,�y&���	c���G%F�A�#	W�S����|�Oگ�. �������9j�C",��]�*�{ch�9�n))U˕�g9 �lpR,�t���*E�%݊&��E���a�8Y����t�,UP�N��]�;`{�O�=I���~�v۱}6֜�v�V�۬�[���1��s�>aϏ&�����A��Ȋ�o�	q�qg�XIO�o�	 �ɨx{�ѽ!D28�y ��3D)U�P2����K[�r�&��ui��^����W�'O�B�űÙ�8SUX��T9^_�O�6-T&������㽌\���r	 �pќ#��r�p>=���4��kr,��o~����I{�'����b#�06����H9O�gq�P!�v]�)��UJ�5�l��	��bpu�[8f�v��O�N�ԯ�����a���\���V�6D��v�|e���@ء�^̋���xx?t�����P�Yv	��}�Oi�������N�'��.��J��KY�Z�U�?��N��w�]�	�B�=��.���jb�kP09`Y�e ����鑊�vSQ����!;��vÍ�И�a�[�Ul~�p���p�eu�'�·*�_�\�
�3�f�͸*��W�B� ~��+_g<�^g��H���4�p,|~c�s�V��3���(��Z�<x�'�����N\���k�����f�zCB\�<+Tq�X��Q &�����9G�>��NT0R�p�Bh[��8��~P�	`�g�ϱ�j,�K����5.�˜��8*�>�y�kȅϯ�����c��-�a�զ�9n�G�m��?f���vɥׄ��u��Zb�z7��"�$ϙ��|7�օ�Ah���}��T\�gc��O�m�k2y6��4/�!K��p%�N�ֺ�r�SI��ݥ��%I2	M��o?=r  �V�5$�*�c�9�ゃ�k����K,�$�L��0&?�0]��2�(Z�����q-���B���"7�o�-a��ڑ�lfS)<�N�QˀXE=#wrP^? �����&���r�J�˱��G8+���� ��=L*��x&;�	�p<�l���\ �de|y��$�ȆH)��\�x�<s 
�gŽ8O�)8y%a�E{T6_ �v�0����617��ע��ƫjJ���C�i�Wp���h<���W�1��1�<��8T�)�8c+uc�x�,�+m�m|��d�L��T%��gB��ӆ!O�u���~��b�l�X�1�O��b�>����w���֨W�~����v��o����R�<���`�~�T@�� ~�y�KV�"���j<4��K��ld|׫M��y��F��#�e�+r��Zµn'�R�s	�!p����v�,����.�k����)�� ��o�ǔ�c�P���cLbb2�$���K�����U��7p����8pЧ?��\^"�(gu�	�,%��v+�;����vϧ?o�yͭ1�O�Ӵ�MC���:�����[��0F,x9������?�X�Ð�X��])�����(%�:��s#LD&(�v ,�ǳи�:
�г���t˼�N�$��㸮T
����C�^q����7��g@�k�l ���o��y1�|/� s��.��`^z��IZ�pO�Oq��2�%�}%Y�_��I��gmb���U�z�}qf��/~�0s�fd/(��u��U�am���S�Q��ԩ/�����=�������T�t+'ӱ��f�oe%�� K�qw�qG�����!)in���{�9I�+{�|đ� o0HA/�S� �1e�W�B���=7I�2@��T�+�%]�*�0���Xc.�i�p�<Q�s��+k\p�E�E���!
�O�!:&�@
7C� 
�]D�4�p��	1F�ǽH�|�7Dq�kHL�V̆��g��'�\�&O- FXDO<f\tVh5�8eN[_�����~�H��s&()��p�^���s�3�OARoh2KO�݅(p�2�
|� 4һ�;���>�d\��(	��) 7��k'5��?�%N^��?�M�`�'����"����K���2
�~�W�\����MB���`L7qc
~Иs��q�0���$$�D!��j=�:O�M�x"�#+��j�yZ�	�0s;AWO4�-# �Fla�y�k_�����7���_��h$��<|$����{���o����iH0���#�y��`n�����ճ�z�W����{G��J���R�8���-���XE�`�����tǄ��Q���&5�V�X<tL�*E�l &�o��oG���^�:���?��k���o�Piw*& )�L��τ�|�.��t�𢳣:��l���"��,�{&9ur��J?��:�/����o4Y']�<Ε�����k  �X%��\�+xC�S�%�{�I4=�-�M%��.�N�~s����w��T	>���@��~kj��W�s}��tw��i�)��kjQ���8E ���&�!�u-�Qu�I94��q�&�st��W�K�K�ubn>����NEIy��;m��h[1x�"�����Q6�'�O�^ �+�XA�"� E��Cf|��К�3���*<�Z�瞽!�k=��Q�^������C�k���@���ђ�p���X�ʅL�ո��K���1=��
~�|�m��tϋ_��o��A;:�����>f��[��.��!#�w+iaxn��p��mb*v����{���Mw�y�i�a�3�r�R��rN*���YC���3����E��G��G�����=�h�c�}"�aM�H=����x�s�
�+�&?�ݑ��Z�i��%�(oȟ�=n�ʵ����@)/���,JUޖ��R�/N,��J�����a�z���^���I�T>�k=�����,X��h�R5��nD�6���U��;��}v�ȂMLZ��C{�S�c�Uצ^���h�;��^��F�����_��CG�J��ɥ�'�B� ���1>��&�ׄ{����o�b����jkN0!�ݩ5vQ�&jUk/�^�'C7s�aW`p����bO��B�iBH��$B�HG�%�R�����ϸ�� ;��� � 2���}�}�*��g`b&kv�ۛ��v�%����1`��Y��8���'^p��][���o�I�*���Ӱ�x�����N�c��ŰW��W��ڤW�J�H,�P`Qz�ܠw��QM��}_�F�߆����v�����1)��u=��k��|��~�-������^m�c��J�i+��9��*���I���DVmrz��Aj��*�5/��~��������q��m�\���P����f>c�Fs`^+i�ThzN��jozӛ"|��}��2.�%T��n$)�5��M	]�ʪ�,TZ��X��<`�6g�Q�̑)�I�_�.jI���S��4b�2A�β#��t
�I<7��g+w��,ƀ1��Yq�pw�}w�0����-G��܀��D�����Rb[wL�� }��۱#�6�y{x0-�7�<��-�Z醋f}*�AkA���5^I�R
LWg��������T'��vع{���?�Ή��'�mj:K�Z)�֤��b�@�D
�6*OT� ����ƜB�yEj�0:+镘6y�h��+�א���_hp�{t|&��C�F6�iH��j/� ��l�F�L�ð�J=Ile�؉����DW��Y�pź�@��)b���$���x8Oj����%DN;6ޡ��쑇�N��Ѱv�Px�m����ID]���Jv��nu܆���~��l�=[��z	�p���ѣ���=�����*�n��F:�险 IS����K���"y�H�º7b=���+jL_�G��C�k�pˀ/x!5��aĠ'�D��M�eWP�*�,��̛&�%�n
Lv�P���N��ɸ��������4K3X�(S��qH�|Fe��d�fgH�++�z�w��Q1���g�$B`��J���Ur<�B����lM�7�}��k�a�MTÎ����I3�N���eJ�c��X�z�σlэN�A�l�L�6�@{z��������]�G�o��]`�]���%_>���zLeI>a��T#RN�fP
(Y|/?ie��3�AZ��Y��>��0�'=��G��s��K������S�k��hRD�7���+� ��EQ;R_x_\����^~� ��IB�) �?��?���>�яFu�9�3p�8��.���Mo��`f�q��ܿhS;-��lf�|�zb�3a� �M��i+(m4H=\<�67h����nVA���ٰ~�n��Ԍu��ӭL�x��>N��f��J����XC�h���Ry����3:]�{Yìk�<X>��OE��t�rS�a�����e8�1+H���}B~�5ہq��ڃp��q��[7�F1B�R|\6����Y\ ���y�\A��c{�SH�p+y����z�1�@[ ��N+� {p�|��d �f �2b�Bh�p�.�ռ�\��a�;bm�����\?���ؠg7��\�
k(H�ݬ���d��S���歜�����vn�f�o�7��pl�q��rC������;�c��^��UKF}T������䋷A�;�D�3�	�꣇-�R)|^���J�Y���_�L��Q;Yp��w'����+������z�������=��w�;�K_�R{���B�ey�h��So�;�D���$:jIe��{�b,@��'73��#ùS6�诺�q��қ�Rܰo����mг��:���4�`Ǐ��v�F-s��t�T �ik^�%7<�v��8�i���j�u�}�=k��W��r;`��B
�Cc>^Q>�V���E�D�*I[�
k�y���}��T�]-W�n�j����	�y]�#��V;A�6�w��."���h�"����9�o�v-�E���+�J~����?��N��R�U��ꂼ�dR
��> ��ІFhx��l�&'6�wz����-;xpq]�����'��z�S�ݍz� ���Ӧ�mo{���c���I���Z,��l�lz�Lkf�Ըa%�'��T�eyT�
C�o�u"����3�>�$jSHҲ�	�A���w�ԧ�QT:S��@���D�:I��D�Aة#�IT��J�ȳ�y6�GwIE�� �+6���?�{|������y���}�I��
����$����f�mE�h�j2�w6�9۶���0/)����I�C��½&��J2��RF9=<��
1��J�$�J��g�����S�7�'6h�i��N�Bnz�@$��V'���k���g��/<C�1ĵZU{|�U&f������z�b�F�T�6vDӱ���Cs ����f����������/^c�S�#q��-˭<#8߫E�6�^ .�֟v�̱.qW��y���'�H�Ġ��^�je��8"Kv�
�KΉ:٣O�%��Q����X}�+���s W>+K�t5R���!:#`�w��X��F/��"��8�Z�G�_.��L��#����]x��v�M/�͛C��cG�
�KF�0q�R�3�� ��<n��9o��mp�]��'.bra&�c�R�@6 x��i*��;�T�3�1�J˶l��c'��?�����+��Ѷ���`��-�N[y*����n�lO;mG\D�¬��y���ڽ���ɵM���`��d�)Xs>�]�
��L*<���'�e��e0�Y�$O�ߍZ�Ռ�xN�UNcxa�"�~��N�Z�}AVS��а'�Tt�D����1��j�XDՀ:]��#�b�0a������薆h0)q����.�Ї>sI�d<\��[����8�سx\7|�e�t��G?�����7����s�ґX#�رV>Lr�
��˃����76�c�q`d�/�`�qL �q$��mг�2Õſjd��������~�ؓ���W�������R
@�Uo��a�#7�l��������7�9d�(�>p_#�Ǒ���D�:�%%Q���8c�8�R�zݰ�Q�(>�s� �rM/�gx��:�j�Z�]�3@(ƥ� 湏�m^|Af ܇���H���dm��ݞ�:;~~������H�z��*�΀������_�r�.�|�!���@Qe^��-ڎ��؁}���){�˯��\zA��ь��F�����
g���p�
���:�Z�X*�����J��#@�C�E�|�7h�~���`�K�G��0�N��'���}�{�lv���P<���Z��zc>O�s6x��|H��k��62kw����R�]|�����-�t 1O1�Д'VH�7�+Me1�;8'M� ^Z*i�h���#hI�tC���F�ވ�����Ύ�,��*�*��C���w ��?��_(���J� �<j���/�F9v>���^�̫2�y�4�_��6w��Ϻ:؈���'��l��4��G�%y}�n:�М�!���f�9}�}�} 6}#��6�ڠg%�[J�i��k������m��>�P�yr&`C3p���pV)i���a}0�J��}��G׶V+� w�_%��^SPG���I�4��aV�I��UN���7��0�!�s���+>�Ւ����r�i��t�h-�U+U�(n��&{�UW�J��2���]�݄���p���۫���>��A ��j�](�������$�����I��]aמ��tI)j�;�o�2l�ਢ�s���K=1���sx.��=+�u���Xk.�/ʕĦ��A�<߾�бhWR� �S!X'F�Yw�+�ֲ�Z��r1�E�)g�`>�L�I0j��)Ҁ:�"��{P���8��a�9B��lujvr
�%9a.i�N��I;>�E�5��c��j����HUdP�T7L��n�q
C���|�)= �M���n�\Vy�RL�A�Ӌ����z��J���ѧ�~��]�v�o�˟^l��#sV%�`���k<&��{��MP1�|�
��J��A�l$8�t��r5����t�xo��F{��O��G��l���c�@��ԗi2���jL��QM���y�Y+W]uU/�?��)��d��mF�W1�
�� X�u�W��b`� b�}�.��Ҫ�Q�t���Z�10�1@|���X���5���)��p� 0�p��Q���������NBf�.��}�ԓRT��D�Und��>9U������9gO�UW�g'�"�[�N�����@�j���?ʋ�9~���S2δ_~����.j�LS&�����Z���m�4k�]w�]�ޫ���+��18��LF>}��k\0 
SsG�%�W�<��4�~R���p��L��t��ž��RQp-�
�J	g���>�ǹ���#��+������f1���Pi,�b���Wg ~���j��-�������㚨-H�9SUd՗�o�_��/��m"�`A����j׽�;����N�s'�����7�3 p��FE�� �H�{"��HH.6���£���T+�x��a�7虢��f��5���Vg�R�f��b���>g�ݶy�:Lj�,9)Jq�v"x+D�x}H���d� ���+12
ʐ���WN5��H��6����\e�P����7����S=MW����c�[�� (�c���L��>��z�Ii�=��tU�ŗR	3ދ��<���&�7�#�Xd7Mc1�>�&�K�i�Ҥݲ��ħ��� *��ih��{U�b�!|�ѡo�=[)�}�lwb�j@\��}��
�;1����f��)]�l�rukTE���h̋�[�ը>T)4�-~A�]T�Hă.��u,�[��:xCls�F��0;0���	�� �F�p>�y��=�*m�g�(S�F�(�OI}xG�r2����a�ޱ���y�,�U�6՘=���h�����vp�!�P�
�]�|ʞz�m���I�:c�&
�JqStPlT>e�j�A<x�	�VLH�td�6�YEi)���*�Arl��C���|���g��VZ���g�i�]w��>�b���	�\�ienm�{婴n�qz��Tд�-�I�trV��NO� f�X�A��?����TWk�[Z'��Ϝ��I��48P}�-6\��AyAh�9:��~�Q{�����.�����'�SOcF�Vc1�HFϵu�i�,%�zE={nj�Oe	��>���#�A��*����X,!�A�l���mƥ�5��۠�C�
�����}�o��O��B��n+��ö{����Q�s��:�vO.J��@q��cJR���{H���[#�9�^'�(��D�LAn�(���@�Z��G�)��8`�
����O8���1	��� mҶ�R��� ��N\��.�#���&��q"�X@[U2'>�
ߠz6SVA���$-���CZX���� [f*<�p,?\Ӓdb �Đu:�k[�ֽ�0je^�w^Z�I-*�$���b=�y�X��U��tu��OY'�5��)�2Р����uvyNЋ��|uoo������rG��V_<'����hյZ�w��B�~�Ⱦp,���#Mb�����$��?�+©�'j�zUF��;@z�6�YI��j\X�额q�Vۺ�b��ޚ�s��]v�U����p�R?�"	��Մ������5���$�� AN1j��O���H6]���Tii?a�DH��Zn~ ����V�(h�!XMt��z��v�^�<���޳c6�W_n��-�Ś�j���?|������ر� {)��HO���"�̠rV�5� ڢ����}�7h���T�%��`�mˌ����[n}~`[�a=um��67_�a�Ie&�#N��)=%�����n7�}J\�d�Mѷ����ٽ*B@*ψ�qN *�Yb�|�Ȩ5_���	���#E��:?D�{Pw��� �kt�?z ����s��f�!�e�v������	�N,�Ƈ&M���U��N�/<��\$�`%����ʡ�ngbX���Ǫ�N����x��2ܩ���U�^?��\��jh9��Y��^�u�l�F&�X�`��;��3�w�Xu#m����v�pÚ��=�$>�oV_��,P�aD�K�A��t˒֚����^Y�y5�O
�ϕ﫶g���ѫcAx���C��s�A�+���*�E]Bw�XuZ�Zu�lG9B�+� ����3�]&�U��a�p�jK�d�)�C���m�����+���w�����|�}�O�(�@���rf�����%t2B��B�op�0¦^-�:��I��l�\��˗_�o�*��Q��4��R��R�Y)h��~Jr%��,�۵!�o]�x�R�O${MT�q �g�}N����=ީ�NY���$���nB3˨ۺa�����R;���?����z�.��j۱����5�;rׯ�t��Y�~>a��A�+I���F�x_d����g�<�mO�XOb*{�D��I��ז���XPH�ة~��Y�/�?9xP�}U��X03�Ȫ�N�����rq���\�R7x_[��	臹wr��}�l�鿱���y���+���6=���漕p*��=�W)�}�y%( "@ݿݍ.p��K(�fc��}�y��(�m�O�4�7��Jm��/��;�����c~���,^��k�_c�-�1Cޤ�ڻ�~�ܯ˓�4�O},~�w�G6������W��N�ju"���G��fX�����o���g�]��b;��K��8����X��{���4�Q{b��=0|<��yU�O/�lW�>@��N�my#�h6�F��=7�XHe��j����@����6-�Vd�S�s�
x�,H���ي�-�O�V��(��|�-Λ�����|�^�����ZDZ-�]^��r5F�� ����Z������-�]�{F�|𵨓��pN��o)�Q *p%�����n���9C�4NF'��QB� ��Ԭ��KI|��+�&Jm�s��j�� ���u�sk��F�@x-�%L1=��LZ��i����'?g�~h���E��isI#\)e�M�D������ƶ��n�����o._�] -����yK6�`+�� ܩ�}l,�`)�����ʸP*���`�����a�^Oʥ��2p)�Z��T�c��I��`��*�D-�5�f��܍��\Wk-8�n���y{��OU�uߗ�|Ggx�2��D%0\ts��ߋ�e����w��'����ˌ��7�4�t�t����`��`F����n������Y#%]��t��z� ����D�2y���*�Ν�2����TT$�U+i]��˕ؿ$5K�6Ab�̅/�%����e17Mx���>�J;f���K�r�C�j�+&	ދ���jSM��_���H ��D���-u�z(��6��v��/�ZKlb�j;��bg��۪�vb�8��.8i�9cX�DuD7^�T=JK`��h�\o�r~��p%�㊟ך�{ݜcNY����a�e�Q�l��C��1�x�t	�xO7<��a :f܊�LO��rX#1�	�-*U"`x#w�_�gG���{��X�e�ڭ�u�i���b�F�Ϭ&Ղ|��LNs��KI#�r� g`!�TCT��ҝ���V���?ߊxLǈ������^W\qE�
#O��z�.D������ܞt�Өݍ�a�������'�r{r-�Y����2����Qi��C{������7��]x���X��C��7��K���:Ҥ�c&ʎ��wm� O�!��:��2����NR���.�kb�������� 5I����r��uXZ�b��ü$L�C�_��?�jfړ�FQ��=���_m��/9��^�Z�
�Нw�Ҿ��'챽Ǭޘ�fk޺j����Qc��h��<�Iֶa�z�O0XA`��H��0��
�k�'���A����7]�.�0Z���Du��k�F�J�lg�}v ��ǜ��*�' F%J��).�)L�)�C��Т�1��n��6�����x�w��gϞ���/y�/G�6�j�	��㜤� )Oe�~�m���.;�^��Kl��h�Fh��l��1=/a�|cґ�G����M���G�~Q�Nu��2����+����'+�(/n��A*3$�z�68鰓X���9ߓAx3Nt�3���#(�,
mPK,�6����a�fw����Z��d��"�i�����(id�ն=�ϱ_������7	��lۼ�fǏ�#��k+V�Xb�����P$�*�DMb��.�,F�RH��ɚ+}�c�@���7p
�����$ot��"���0�SS�5VGt:\� ��v�M7�ƞ�Gkr"(!��o*�;�������P5��ߒ�g��뮻b"旼�%��W�"ޗ�R�q��b��~�R��,�O����-��^�[��T���F�h|}9\r���,�c)Z���~�䋤c�b�l���A�������-����v*���>��������Wx]�w���뢟n�����̆y��,� i��(z_�( 0^bj�wۻ�h�O�$'��1�O�Լ��� 9���P¨T�F�w��ٳ9zE|��='���/'�ru��@Y	x�/8B�0$v��/}�KG��e[�� ����_p˔bS Z�ت��涬`��q�0����m�{�����}�=��S���J�̐��ΰ�$աc�(�Q?N:��P���J"�s�=�^���/�rs��2���>�у<!�d{����)�ͻ�~9�V��f�R�ӴV˔�?|�)+_W��Zf��"~�x<0D���6�1/E7mǪ%���K�r_�Iu~�si�K���dƻ~�`�+�8�����t`��~��n��Г$���uJ��-ñ<��#�L���g�G�17�s�OJH����~T�W9��4b��Rq�T׷�h��G��"}2��)�I�[���Cf׬�J�����w�"�|�gon$݁y���3,1l?��'��R`&Y&#��V'�jWVs���;��*a,��G����0�m'����l�D˶��;������<RD+���^�M��z�z�9\)�õ�R79��L���J]�q�6)@ə��ԗ#:�{�qn��U�P�8f՞��X�����ʓW���fl���:��`ɔ[���a{�5W�A ��x��hx��I@'}.`�\��܋_��8����IKW��?�S?��cء0 ���cy0��a�<��|�3C�/�wa�,����w�=����c&����2���aB#� ���{�>a����G~z|�R���Y��1��8�(P��n4��� �Q�
��`���{@8U��r�23���/��[� u��Ja2�ݜ�qaR3�}�n��e�}!��ϯ:�=h�ő�d����'$��t�'���Y�U	�>�po��N}���ə��ONTs	�q�����Tع$*�$jb���[:�|�[��{�id��)�r��$΅X��m}?��	�pȾ���>���h8����;ڶ�:�\{�tû/)=+ 2�06���	�.��(�mw�����k��Q5F�+��2�� 0�l���1Q���Nػ�o���3��y�e[o�˽��^���[qΈ����ΞC�Mn��WLȭ����~$}�~�;*�����q�u���9�~~:�Evm�nZ���ޭ��׉zǩ��x�7�Y��?�A/���׽n�v�����K�
?�^�8�Z`ﭷ�:탹9o`��cp>�{ؐ���
7�|s��*8�O,{�XjG���� ��r3Pzn�|�}~CJ����w\|�nL,�������7�G�%��q�q���"`�2ep���g�Y3��!�9��J��o���1	=����~f��M2WT���J��q6<p�C鯾�t���:�6v�����P��l.�n�A7�[k)[�[7QF���8�=]�p����h����r��zʠUp߭\���y�G��zg��b
S{l:�L��섃�g&���ի��,�O�1}��ۋ�@����u�r��9��m����"5�0;n�`�m��n��c���aTY�)}���D��kw�-����&[l� ����T��׋ 9�4�7��w��&���5��0 �[o��m�\��6�ݥtp�ĵ(ӃS���F7=`����ݕ�3wB���X�N�d�J��Zݏ�M�� 7`����������;�i�F�"�Hl���z9,���T.	��>���旁p �9&����Q�;�nq������4����@t�w��/D�$�(�iYII}f��er^���"]e��`~PU1���y����|B�LRC�h���kl�	'�
d�,�
0�c�-�&���Ғ;HKt����u����v������ݻ���t�=/^9�m�	g�h2]ty�����t�iAZL"o������̛�*W `��g^��l�) w7gyj�/�NR�*�<��@��P��T��!3D~�F�ϚBv`j�޺�1Q1P5P%>�&Xiky��"==VǚŊ�?��פ)2���e.�.=
gBh��X�2UҔkPڽ�NS�?�$?+�^DƵ�z�����u]Ϝ���@|� �VZ��=�I��2�k{i�����d�ʢ��]ߠEX�]#:�׌���*��\r��bV�̒`Ɵ�ɟx9X
����o�?��OA���� ��� 6�͑Z���'hͩ�3�������F{��Z�n+��S�+ƝZ��ˢ1�㼳�q���4D�q���(�VC����x�)�iB�c���(�x�����L�W\�R��ot�,���<Nn�Ml͠����F�&Mz.n��0�|v:�HJ����:�w�r1�k:"D���@7;���C���ܸ����x4q�Y6_g~e�L-:)�a�c�Y��ô�������eS��T�t��j�8�ndǇ��d�� �=��)𬨦P�h�v0��ݛ��o��t���7�������0�qݜ�6\E����X5N����6�������^mV���TL�S�M@�aX�g��J����4��4[+#��Cs)R�eb�k�ήk�B�6�� �:�u���O�{��g�p��X�Re�0F�$��5�\N6kM�r!{ՅM�?���1C�5���x�);��x;e�h�9.���bn�k��֣�!O{2r5~R��f�T�Kf�h놌�C"�����%X�i�$7�$e���&`��,��g0�^{�4u	6~C�����+L�`��` �t��m�:��al��Z�r2��Fo��G�������j5L@�$���ÃE��]�yԱ)p�=��WC�ѝO']Q�0�����`g`�"?`�f�[wh�_۠��R�/��Yh��d7�7��)��� �ڌW�U�&<aM7%(ޘl�&-���U����	�%�w��`Ǌ/f*W�'��@a@�!��+;(�
�^#cR��D`'�\���y��I�Z��ʺI~�2���r!����*���SG�y(_1��?�����o��-�T����y�SGdfХg+r�9('��9󩗳#�	sϵ,-7�l�����^�� �XTה�C��`q� l�L8_C��,�&�ՙe�u%h`e��05��Ɠ\�&����q����&���Ν�Ƭ7�wҀb�_z�F���(�!�Yk���E��/�y ��d:�S��׌�,�M߃�|/U1�ħB��^��ċ�T�Mv1���������X@@��x�K_�{���Nf�	��Wjة{��>jU�~�4 ����f]�E$\�i aDv3d&��sB�$�`�Y1/GuB7���L�z��1-�E6>�'��I��?���/��/�Q�����漊���G���ƄMjV�M��M=F�0v�YXX�L96X���&u�Ė��s�i�S���ߑ	ov�0��]��ls�曞좲�Q��zn�Rf���-:�ڰ�ONIU"���F��0j;��Rׁӯ�0iR�9�7V�:C7�R�Ә�w�^70�pV�{9��N�(;�r��4�����{���^���:�(�iH�s�� U�
�E��`�M� �|Î����V��ͅ�7i"�f4�;�j`�,�,g���,��<S��l[,-�=@��ݘ�h��g7v���|e��'��j��>&����h�NV4�ko��38�βobc.��q���zӨrF\����`ves_u����m�ct��p�MZ�K�A,?E���ϵ%4�����k���{DǍf�F���w���h��3s�����?O�*C�t< �m�N�U}+c1���fl\NS��q�{] \�#��S�z���*[Tl2r���r!Q:�dZPؚ�KD�����U���~�{�s	H��7���Ƙ%86 ���񌎘�9b�p��G;��!���3;�\-��C��iV�`V�=�W�t�y��w�!�`b��k�R���s�Ygo�EY90M�{Ӿ��^�*7�tӷ���t� �y�c.H^t��ڄ����ܕ����w�K�R�������=�
��t�y;�y{v�]����8�ԛB�`�n�)�{�����t`ߡ����vl�k��Ҏ��}�:3��B,AG��rz�����ޞ��=�q��V��9��L�^r���p&�H�)��BsF=���Vc!{�:�9;ܹc)]u�S��h��Y�ày���r����ӏn����ђz��+.K�G��j�QҘ�"�{�k�������<����5��\�']r�cz���MtG�M���O����v�����a����.��ϑ���ݬQT1���V�������}����;۷��'^�ce��j�*�ܾ3�|]�s����[��H�:5D��ID�����[�n�N�',gg�g����{����$&�:�C�ػ19ֳ}�N�\��I���1I���Xh��������+.�Z8#ӧ�a���}z]�|�h~�[�?�=��v�m�m�3vs�� ���MjB���AP�� e��Q^���s�Hm�B�򖷤?��?���w��镯|�w��H͓�Dq��(��у��o���FI��ǋa�J�[����E�xvO3��qV�j�*5�$�9��$�5���`���7�"=�9?al���*ؿ��vdlhh�뎝+&��������?�A��m ��=�)����
�L'��Pڶ��:u�E��qR�x)������ޟ����r�������}B���~K:��mv�5��^�Nfs�%����t�?H��;�o*Lc0�u������ғ�|L�/vlْZ��Y+OVӶ���߹#����?��H�{�X��_v}z�k^h�q6�:���n������O����L+X�k��	�����v�*���t�u'��c�q��*>�_|��?���j ` 5�ϯ�ӿ���O?��K��u _���<��csxם��o���j��v�];�W^����/{zZږu�uX�v�D
��߳绔�������7��Z����7���ڕk(8�� [[?���qpUv��y�_���]���²}!����o���9m`�5[��m��5���(�/~�o����-�y�^�����;�fK�s��.t���瞫R��ۇ�_���TW��yn�L�7M�ұ�l�i����d���կv'k�+�FK�L2�@9�d*Qx-B�ގmM5f�Js��������@�@ �����).�S��uf����ɍ���t���Ä�Fe�0Ĉ���E�A��ʰ��7�t�O2C:���⃉Ԑ�W,;���#�!�����[3�ܮ���{�8�y�##g(~�c� =�����Y����t衽�k����M���1�]|ۙ��:Bǘ��`�}֊��e��iea�30:�P8{q�L�V�껲��+7���g��{��ťIZƙ1�a��@���R/8xwN��Xp�_Z�Z�6>ҋ.ܕο`[Z\�}���gυi߾�n/�+�}�bڿo�m�����$j瞳�X�Yimx���L�+;L���}G�l���x����s�MȏL�䒦��/�s�X����<ώ�fﭥm��2�ٰcV�%w^��s_ ֖��=�3��ڈE�w�z:��rmt8u!�Hq�&�� �m5���`Q������Ε�K�;w���&������G�`���ׇ������w��cǢ�k*����{�=���\��=hb���d��c�K�&8V�wl%؏����w���0mhl���Ǚ��si)�d��k"��57'�Μ���2G;�1k���dSM֎"	�j���s?�s����8_�?��F)��Ϊh
%y�E|_Z��R�-X@M�2g�8��j���h���wZ>�i�Eg\�L���.��0�
fw�u�1��א��pF� ��rSq(>��F��D��]�z�� ,Db�9���w��_��4K2غ\�X�Ԑ�@b�ǉ]G�F,p^ٱ����4X\p���]{�=�ܛ���Ϧ���<|�IO~\��T�ڝBkn/���7�wpݓN0#,���T��|�[���HKۗ�EoOW^uYڱۘ�;kvHM`;]��J���T`|�onM?�����祧=�t��%�\�9Č���QV�D�����Ӿ���}S��������fl�{nK���µ~���� V���i���ih�S7|5�r��5�S��.�e�ԫ�'nӦL"���@�+t0؞�����w��}[/���������v}�=�^�Z��YY�vC��m-���;�}�>����uO�:]xɹn*@��:i?�����:;�*ZZ���7nN��v�k?qՅ�k���pSHi��2��",Uǳ���Nnڿ�7�J7~�oS׮钋/HW_uiZ��w|���&� 4�b���?���a�f�������A��>��?�t�y;�ֽ��y��Y��<T�eS��L�uwJrM'[�d�!b�)l0�}���;  �$e���ou�x�^g��������<զ�m}�(㖡��vk�I@Dx�v��=F�7�҉�[���舜*�Y2���w�c�w�d�r�25p�y�v7C�(���Ka��FdV�YV�����X�DH�Ƭ�A�N>yI���P���*��"�b�����,�}`�1�>ے�*<����=���ƺ�����ϸ:������{�Ys�0@XXr��`���rE9�y(�G>�����t�w�sU��O>+������W�pj�d�f堟��J������o�f���{[��M?0��۞^������Zc���3]J�Rv9��D�Ů}�a��?�����|��I�Ȼ�yOO��S�s�n�Kf�\�R8��������������L�?K�ݷ��ql |iz�~%��ϼ8��Y�z��׺�I�(�L�կ}#������������Q���_���o��0�N��~�f��xT6!][/��[��O�����X&�~�^�^��Wÿ �&�lnM�3�<"���q�������|6����M{|�M�}���[��7�s�s�	%;s7��ܷaZ
� t!撾��/���_ߖ�}��3YL�9'���_�~��ޅö�g�~���X�6[�ϭ�ݟ��~{�䧿��eb�����_}ëҥ�{�=��L��n�� ��l�;�\��/��j�F'?"���l�z�����Nn�U�H�����D!m�������l6�p��}9�-�Z��3p~�*�5Z>���mm�}�<L)�j�i/~�En(?� 3����R�)+�4�a\��&��ᆙA�Y��|�C4�¼�ı�I!�ɟ��������n��
2��Um ܊��9Fu�̈��m�,���ݾ���s�1��N�}������ie��tۭ&�׾��t������jKS;��Fͥ� 	�1����}���M������|���L�_��t���9�r��]��.�[�X�>��/�>�۟Ɗ�b���}0H�x��M|��Ya��	�*nO�z�uS���nL��vȄÂ-�s��>����g~#��k^a,|��q�s��hB=�ή��o�bZ��������a��ᓷ�]g>]���`.9�Ф*ܴ��Z#������_�n�X[pG�n9����䟦�_v�;��3��L@.��u�'>���?�t�@�7X�̯?~���%�=1����gɜ��s�Y93�&ﬤ[~x_z�{?����E깣���t_z��h���ڼo�=A'��,8�h�Z@��u2}�+w��i}������K�Y�??�쬍���������7��`��JkƦo��W�ܟqM-�h�?��Ϥk�{F��1O�}�͝��f���3�:�&,��)�O;A�v^�5��[���o@�=+|��/ RMt��p�?��ϟ1�g	^Q���"ܐ}YF� �F ���O�[��F���َ2L�K+���w=���ȷ���/В�M6��cp3$[���H3=I$�M06�����G?�Q�j 3�;��_�r��}=	�@�H��I�A2VU:�!��Vs�=x�����T�r�	�����z�(zg�mw����~�Ύt�}�|���~�m�o{� x�c�z`-=��aS��H/~ɥ�{\�����c܇:���0=�qW��.�A:��!b����t�}�l��I/�k���.cav��('X�]w�7 YN�\�Tcaw{����ko��>��]隧</]{��y��84��P�m���xMZ?|K"�r��NS�/J���~��������[��_���-=���٦��KLwl����-y�k��ք�!�0پ�"�d�Ԙ�iI��, �k5�}h���K��ړ�x��{�y_|�9i��a�׮����_n >rf� ߷apv�ѭl�[ץ[{w�ZX^��`���M�S�v}z��c���y�����G0ƾ�.{���os{��2]asp�	�U�OI/{�N[{�j݄����Qz�������Y��'<)=��m���*�g":���g���j,���RK���w��Ɩ�t��ķoK�{����9w̕M���m��~� |��!�2f�i�9
ႍ����'?ُ�}^����U8+�Dż���o|cZF��������	����:�`��{�= ��`m���D���iˍ3�'C���R�}�.�8�\�X�*֝7���	��H,J�1�0gl=H���8���JkH4��g�� ˎ�0�hw�)C������8�$r� �
MS�����y�����_�m�/��I�7�*o��u����)�f���$�c�Է{^Z�Ą!y�}gүy�y$l��6�!�xki۲���*=���LO���.��xW(����ܟ|I�'/4�u���.�n0�=���%D����e\�F��^}�3|V�����H{ο��m�1�����Cv���HYIW_�ܴ���;�{�%��/6�Z�ݻ.N�{�����Ҡ;p��ֆ��+�N������v��f��"c�}�����r��@���u����⍴z���򫍑ߞ��w?�g���>���i���t����=+�֧�&d�<P���g�8�oH��zz�ŏI������� ���_~��ߡtnS%�X`>���Dx哯J���-����<-\c������'�N��T^�P�8/p�l�����g��o��w.���g��;�\uͳ��������6pX.�����级>���_�YyT~k������0ը!�0�#��+��}�2(����I�H@�d��s��9��h8�L����a:w��UD��}���������@(F<�D �+;��g=��6���"8
E�5n��g�
&�����d���.��ff�X�Wǅ�������v4sB�l� ԱNv�J̋��^�Nھ��OT�"Z�ӵ�ޖ.X����O	F�I�=�H�];�2}�C�P/K�lm{eg��Q{M������3U߫XFUM���6u�0-�c4,�Jc�;���o�(������ٿ9*킁ނ�gl�ۖWҶ�(���z��⒛P�Fa�E?���"a�Z�<-~y����bJj�d�K��F���a���:��AG�3�����+9�7�ذhs3�cO�q�� �ޘ��E�@t�r���X �Ѹ�����\n;ǎS�5M��������ߎthx��υ�<#*k�vb&|�&��\^X���HR��wβ���!*�fI��{6�6�E�ڗ0u��z���p��g7��j��/,�i��0H����ǀ��	��D0c���i2J���f�q4�'�/�Kc>�7��f�JS�lDՍPsU8GЖ!��髮��q�^B@ ,�p����O|�΂�5!x����c(�3�p�IB�.�c�2�����B�I�P�Vu���#sC�����%7Ex"Bc��#
�5����F�t����sD�{, �� �08�U�v�D�t��*�]�G���މ{��ȹDכ'�g	g�VX��.j2��6q�==��3���Ң����7�j�Q�x�3�6F��p��M���9
Ï��f����
����g7L�+��լ�z�_� �v[��67y�02b>�3#�k�G�NuN
���^���4-�H*�q�l�.�q
/5J�� �g�"�n3'-P��.���Ǿi�e��+@{�5<:��ϻ?O�i4��s!�_\1�p���� >���Z��3�e9���mv���|�x�:������{L{vc��2���Mx�z^��0�%7I!	��� Б�6XH�W�=�sm�p.�^�Jj*�?���I�	oZ�[�#�b�c|��͆$ŐW�m,5b�#���/8�&�S*�G�:Ų��=G�l�_��צ�'D4Ci�¾W���FŨ;���7�JE�}��^��-��0 S���L7�B�Q��6�P&��u2g(��RL^&�'5G��r̓���[�f���L��@Ք�TA�"���ey��\^s��Y=���&��7��sX�d%Ϥ#���d�qΞ�S�F�I��$�.�!y߰�S{!�ը{���+]]��R���L���U��笻^g��j.%9H
��f�E!��Ef�9�?98�zJcAU.��Q����]6��P�zmfϹ�p��� �N��M"Y��P�&��g�7g��q�\gѴ|ϥ�X��x\n���{��)�#B�:O�����:.ܜ$�Ru<>2���g�t-)F>�0��W�x�)��r[�[zd�t�"G1�U�u!��a�؇a��F��D\�Xs<H���`�0f�UL{�uaNf+B�8畣�M�n��N�iʏ��V��*�b��t�wѝM��8�m������K�P҇$#�JI�h�9�!G�	ozϙU�+���:);_:��C���R��%|�k=�^���T��=���uP$�"��!�Cf쀵�NYR����E�i鵅�^��KF&����L�t[��s���n��5*���-s�aS��;]Pns�j���)�$|�^B�r�aO�����'XpG�g5� *z���{�lm��IE�β� � �e:����R2�:ɵu.���z.VD&X��5�&�'�v���GUj�=��hrHk	{<�Wk�i��n^�Qo�4ʢj�q!�M�CNZ��Ir%�f.��I���M��>��p����h �n�
@-׻��0�#{�.4";�N�oI	�x�D�M �֬���1q�""���QvGͽ��l�)����"H.�2�4dL�$��r@�ט�[��0!;���R�o��T����#���2���C3`i")S�i���)��M�t��u״�:����sű�5�Nw��~Y�e"�k��s<qSϠ <+�i&��穩C��y�������۰�:; �IngT�3����=���f]%r�G_c^S�x��47��*�����,CBB��r��=sM.�����(�.��Y�tfdE��6�Ԕ���$�Y�^�jf��M)�
g�.�oM� �� ��2w���E:�Ng<7��2�\���	����!�^
�!^��>�4��dVߝڀg�Xv�G6#��lLcDS�!���Mْ1+f�>1<3D�S��Ĭ������r��*�̖9{M�mU���@���p�Fs��#�jK�n�@�����~�dU����=C�EaX����j��+�h�6��eS7b�����N&7��VPPʑ�C�̒�q�4Rĕ���}�r��\X��ISƱce����*���2�z�9/�6<��Cv�?�l�g��F'��>�s
��$�G6���#�g@S!rŃS��Ռu��V^�`2]�̛�O�z'g���Q�l�.<����KN�0��"C���^��9Fn2��{^�$g��ba*�>q��J�Q�g~�n�/ZC���$W�΍�C�GwT5�N=[*����ts͸)�T:㧤e��k�*MKw֏l fDBv$��~-�[<�2��%���������C;�k�i����`g^�ٍ����p���^������n�*�#�{a�5)LD�� ��0"�̈봰H��<�=/�΂�$�aE���q�e��Ȍԝ��ȩҶ���=Kk
�tHn�$�  ��v�\wOz�o�d�����>Eo���X�d X��r���r�m�y��>F��g�ts��<8IdP���۵�^�-<��	�����٨���B���Y8"ȸ�ŉxo@��Q1�M��XgR��}�����$C���:^"?���gsI؞/{?ޤv��3|�˜�[,�B/���M" �t���\��>��T��Ft����\E��M���~t�ML���7lf�tt�y�8�7�m!u˦��x�S���\5fi.��1�{HGf4�0�]Y	�cz	��n��9���.�Hɶ��7�@PW5�u��,m����VC�y��C�4�����HGd��>��[o�^���ﲍ��,�w��^�|��hG�1P�g2^M��Fڷ�J_��_��ݹ�q��gv�u��-`�ݎW�"��`�5c���ލ�o����`��)wi��<�t[���Kw�������������/~m�T3�k=s֥��͂&r&���<c�;߾՘���!egdٰ�ƖI���r�GUӕ�������r��D�2i &g�i?t���3�MXw�q[��WK����gբ��ah܃W�릛o�݅٨��B�*W�-9h���D7�l��6ގG������ʴ����}�f/���V΀�ٴ��g�
�1�Y(r'�J� ��fW�ą%C��n$�C�	9��7�!{w򵔷�#���i����XA�N,�m$w�͔>�ZβK�o��7�?�#��B���'�Kr��S�1���Q�ěUL��l�
Q򇘵� ��$][m���ǅ���ŏ ����r�ވӀb89�=��m'X��7��8�}��Й���O��~�L�W�{熬�e�z8ruvu�PZ\�xA����� ��>�ZԒ@ƌ�{�e���}���l﷍��[nI��r[�� �9�P�N�A�����%�O}�=�>���h.�C�����Pbp����v[q�{�M\{�A���#/0��b�������?8:��uS@��e1[�5A)OB�;��d��羐r����jb2�%�=�Ո}#E��[�F�~:D��M&W�9S��Yh@���w�|��/ _�2@q}�o6{��>�;���Ye۶�Ё���jj�i�K�n��{䐔�FԬ�X����~��x4I��X�!�N�\k�Z0��=':�):b
��4j"8����S��^��ь��{1�WJ�!67Ɯ1�Gژk��K/;Xxo�D0�^�4VQ�;jZ�$w�岀S�sa�!`�c�SjL=>?���z�hS����rn��x8A�ڜ�&9�id:j%M�a�;H����ZK��VL|�uK[���?�O��G���x�[p7�GM���a�p����Mf��z����7V��q5�~{#��z��Ta��\��0�I!_ل�\���jԉ>��oz��٫aj�7n|�e��a��ٳk�Xp)��3ہ�����/ki�ӧ��X��ςU�@pv����LaD���h�Կ������Y��r���5N=�ǽp����QB�"F�Q�{��*���%�b��5?�X��GS��Gp���'�0��������S鞋w���n��l<R`���Ю�|,�,���@�Ld����n���s���]��Un�w{����Z����XSfԜ{��G��4��(����^���Rs������h�ߏ��9 �@�q* �l��XI�A3��b�0#2�v/��1d��w:!�9�ܖ�N���o���jb�Vj�!� �~�匓ж	=���ϑ�2���8���{G����1�9Nd."��w���8��j�ۼ��s,sq,�u�A�I���h�TY\�@Q8 Sf�F�L����`rصK���6��T���U\x���G�>ua�p1�!J�^�7-ƳՐ���+��x���H�=/��h�?@i3�c1�̘��N���@|+A���JA�vm5�5/a8���hю��=H���1Y9��J���#�K�e*���Y��t�h[f�֖)�ũg�ոWl�
~��s,6�;��a J�8�iB�_�x�hr�iYu��;N�p9����X�D۩�՘r��9��\�����^[�c Ȫ'#�nd�1J�CɄ�* �9r�+�͜S��G�r�a߫�x��	�ˍR�Dݔs/s<�іMц�Ր݇�(%P��TH��yl��؝�8&}��'B�[s�Bu2��p����6��.&+��-bHk�DA\����?"w��[�s�#5��L���#���b{��%_�t���qH��a7V#Ou I@��,�*�VC�+7�\}�Y"� ?��0�}���ĉ>��}��sr2��h]��:����k`���53d���8� �*��QR��:7"u�Ȉ	�Ĕ�b�\O����֖ �+=Uc�
h�#s� .%*/��R�LD^��ƹ)�@P[��XR����%k0a��8�{3q���S\��=q�m�':��$p:��cqXI;;U�hL�s��#��4 F5���0���:�I���d�M���#hSϜN:&����$�P5��Ԙ�����ܔ�Ʃ�	�`�����M��L��27(^s�5^(l�$M��q
 �&P6���ƞ
FTV�TS�8U=����z�k_�R��`��_��t����!�>��O�}�C.T��q*�t�c�j�=����od���Þ<�3?n���xQ"�e/{�W;c��Έ���/y�Ko�7g��Q  �B�/������Ee*�v�, ��(�IsO���/SEÈi�q��#�aI���^L��q�k�����E��7��b�X$�@8&PPY�E?�'=�I��Y���4I<�K�xz�=�)OI��|��ԧ���˿�I���y�s�?���(����ʝg�?��������I�u��W��������I�f����1\MQ|����E^C�أ��1������{ ��C.U�2��DK%lm�0ܡ�XJӛ��*��6��=��t�嗻$�,@�_7�D ����(ō�l���`�0�TJ����C����5,�g�a�L�����O'Oi�qB\ęqf<�" b 2&��U�J?��?�c�d ��i��	�!���gz�`uw��{���2Eo�c�; ��=�y��7���M�Ɯ�p=�6�d�N��Ki�6r�
�4h�y������IP�O~�4I#$��!�)� 3�8^��:8c'�6��1 �4}�+^�7�g~�~�M0pu�PP����A~$�93Ό3����){F��`��׿�����>;;�tXva��x!}��캊C��<���y���M|Qh���&�NEQ����sc��pq�wp�FnRࢸH
�sQ2l���xj-��M�LmF���,���V:k��1; �L2��x�~�����Z�r
%�q];3ΌG�P�����}�5�y�)Z1L�����܄�S?�S���!E:�)8��� ,��"*"Q��`�;ǀ$�XD�:��&d�����jR���b� ���L>mo��I� �0]�$�I���x!9��w�N�����i����X�Vc����[aqL.��n�gƙqf<r��%�e	^��pѾ�����zM]�g��$h��`V��g��2-D;/�rNp �[<�A$C�6���	�I]vJc����;��p�!@G�MIރ�"q���'�C *�	R�/�5;1��b���Yc�A�5����s1�?�3?�Cy@�p�p���g�?�X��1[b����L� ����ڵ�?��\	�k2=/yP��l�;�+0G�#ӄZ����t�UQ�+־�&|ʣ#�bSQ#<��[��x�ށ�2�L�)�q�|N���XP�C�d 1�)�c�m�&��_��_w�x��L�G�>��Ϲq�@��Q���V�*p�錝��83�e�h���a����T �������{y���/Т�  ���A�wԵG�l;H��bBS�#�$��WҴ����pܩ��Y�+:N߉��瞻��7����2R���
n�5���q��7ߗTSz"����;���xA�U�.�G)6�����ԣ�<?���)�i�S7�+UD0w������^o�Xo��\������vѣS�-�H}����K�������F_)X@��W���t�7LqQ�E�ٖE ��M�7'ƫ�f�2�x�F���ٻ�'��EK9�q���1�=N���M������~ћ�E��g���ȉ�Y��thW*��A�}��w)DV�7��Mnfrc�e�Ek��g�ԤF�^�;,��i���k��m~;7y̽��鎿_W['S��c>3N瘷�Ol=�e���"K�c�����.7E��oH/zы�������o�qjj�o� ���
]��H�x�j�����6��P��贿�o
�We�Z��Z.�~�u8��skn=T�Ͽ�)-W\�nP��$V�<C��&A��߀,L��~���CJx
���u�sI��3�ڞ��8��3�f#��4�̩�*��i`��������W�ES�*��)�K#�3��8]c��?�<�Io^�d��u��-N���L�����b��a�Ҷcy�؊(�=��4�A��{D"����r�m���-A�c��锹=w���`��x����=�t1\�b�f�����\��4�T�"1d�����=�d��yX8������Όy8��:����y�{�u[�W��zsQ�<�Pc� l�R4t'):�ku�83ΌS?�懶Y�h�y�8��&<�'��w�=&HH�˷���C/x���2?���W����>�'"	��>�a%��=*��\:S>�U�F�_������M)D�-���\��rp2�K5�Q�1s'���*{EG���������&�8��b�����.[N�Zʠ�j��g�
UΤe�\C��(+��f���j��jG��3�Q��B�c^g�����>�>�6T��?��� F�c�P�� :
��_��+���%��MR��b�ص�+p@X�h%��!�Z��g��oxksĠղ]��<eY�]g�L��AZ_��[5�i�t��p�ܐ��	l�HX.�p�v�vM6c�$��%6�	X�R�e� ~,C�Y��1mne2����g�6oB�wJ�0p��:�������b��c>3N߈���f�Gc�G�����T�:`�����w;�3���%4b0 ����5`�� ��Z��`�2/0�a��e9�%�q8.x�5t�3֝����~ԅ^W�l�U+sm`l0O�}uX��^��Û X_Ib�
��
�}�P$1w�,��!;���m�]~�b�T�GP-�m��)��+J�#�i#cq��"K�c����ek
�9�Òs7\�Mg��,���3��3�4��bs�&z4s��z@�}1ѱu*2WE�0;���o87��%��5@�$0�2X~���*���1Ҧ{�]������5d�I�i�\vG��	
�$1��(���?HW����(�zh�n*'^ �j����3��"@��"�H��*!S7H�5�Zbk@� l*+���/v�ü<�R%�;�1uʀ	* �1l&a�*���
o/�tS�-���t3�ٙ��1m�әqf��!�Nb�G�cq�EU^�SU>��p���'{���wyf�.˱j�@Kam�0��`�I�>Eq� ��5���\��s�po��焩�Qi	�rFk`C���|��_N?��t��d�ét��3��S 5�����_���}2e_Aa��+8�G>��h�X 7�:��ɐab��'��>�չ��&[f�t8�,�ic�PZ^��h������x#M0����,E�Y�1����pL��N�tf=��������P�6������S9A��=����L���L�G֦��0�ΜxM��暡g��Bճ[���u*���%�ߏ�i9�֔3&��S�RϺ(6T�QlI����[�T����Q���\߉eY�7y���b�����o�yf�V�<[�}F߈�I���h>�-.��0�;Q]��6�G��BW�����ǵ4o}i�D���*���x���Ҍ��Km�M���	u�͂1� �	+�-�װMS2�h�M�>���2u�NVۛd�`����>������!҉UGX7�E�bPzng���~��n<���zP*���u&���"Rڳ��c�����`�t�[V�k���0{�ũ�����d���R��U����Pw=�Mҳ���	���`9��Ua�f�<|(�y��k4W��m�3��D��6��ɟSP3��kk.cXN;����q��0DE��,"���Q��q�ц(A�s��qbcƨZ�dc�dLT�E0�wb�,�������lϟ%�d��rZ�
i����k$�g?����磹��IQ����9"��ׁ����j�;�u��p���k�5'���	J� S�G���I怈����b06���ߔH�%0)��������	�;h�C��N�8j�e�=U9�����v�^z�S�꓃���r�jE�`q21 0��=��J�j)�Z�)<�X0�I��j������l�?h$�(��I����sv�z����0���4Y7 6��v�^Y��tO�p�KȞ��~z��Ҏ�.rޘ��λ�I��E1sv(�$n�MϠ%��_�U�aH����<��z��Њ��^��o�TF[[Խ�Z�uEO��'Q�n3�M�v[=k�|E�C�MM܌�P�5��ⳬS�[���j�<T�J�V��GdB����D ��� MZQC�@=G�T��U�a�1�I�K�����c$�T�ڶ����h�k�<\l�B>J�ҵpm@59�t�|����<��`Eh@U
S�	������o��?7�#!%�*�V:�q�*j�lc�䅼h�nf�D(�ݻ�A�e)y�Z`L��j ��&H\n��b�I=5ew2e�d��L����������mS�a:�3\�����0m�Hc�i�L�o�;�L��1?$n����z]S��:�ԫ�>�*�Yl��`p=<lm渨�����.��{b~����o/J�#1a͹j��D�>��f��jck��Y�X�|Qx�"Lb�z�\" k=H��њP�n	3�(x,�{�f���	7�Pe�X�@�)Е��c��L	F��ya��9��F�>/� �}VM4|F�s]7�M;ZC�5�sH�E!x2� [�Yb�c߸H�tj��� �-�^aN�_�������7��y�w�|E�TSq��xtsD�)�d�OV��^���Ƃ*�M�t��܄<7s0^-ˈ�$Q�e0	T�GRi��q�yO���g4.�gK��b4d��c2flG6�P0 .�1f�I��ii��a|Ua��h@�En���Y/���{�nV^�s��$�z���,7f������ʓ��`>����N�P��h��L `��uIeBj��GtrD6�g��1�R#�H�&�X5jM�髽�/�f��\Q;�J�om.]s�=��hֶ�1�:�3����Q����ɼ!����(��֠��.^׫=5�v�A\x"㎎>�qt �[_�2��������K�A�F��/ӵ�=�t :�	�C#�<�u�s��^�k��jFDavl�i�>�z�2ؕȎ�v3��Q7��Ҡ���=(?�
*��D��ő��a��E�h3YZ�L���5ǖ=O\�Q��h#/��*��Be�W�lA�vX�^����~�<�*���ʩ�%��Pc-��0e�,<dc��R[���b޸g1Xݣ�����Rs��m����ܺOƑؖ����D{�
�G0��#��Jz֑-���)@����5�_	(��~�di[0�L#�D�b�1����������"���~#co3F���Z,�=�q^%����H�p$տ�^۔��q�g�&2Ui���ccp�cQ9Q�eQ��פg�\D|���N W@�-�����x��=#	�h�kk���p��V��B7,<�A����ͤ?L�����T�B):,Z���iqkB��8��c�6H���&XFcy9gj�_~�1��������
�#T��Sy���T�̀Aẜ4N��ɣ& ��Ttlsv���y�����]6�v�T/چ���0�5�V���5�,@�T��E+�)՜��(�E��&&�+۶Y4*m��Y��)���H�"�^ڂ�k�����F�?F�(
�m�՚��x���<en�YM�X�����^P	 1j�p�f���5q�<j\�b��]ku=Q(�AYj{M귀���6ؗ1��D�� k�k�ه��_p��ڋ���Ks�&��7�)��s��k���#�(��υ=*&K��f��ؽ��Ә@;lʙ�%�WLL�Ɇ���ʪ���V�d��MK����~�Y2����<�ԫ|;e��~�I �669���ML0�k�m \t��r��oRx�v~�H�$J���.a�ndw�m����[�M���juu�Ȝ��	���?7=���{|��Ճ�7�;���cr^g_��������~&��{ -�=%c2��l��;�W�������=�g"n�8X�lr���[F�%������g?�m�b�Qk��]���Cj��72�ig�V%�Mt�I�s<� q�j�6B��vZ�A�^���CmU��(��@0���2ma�� ��ԧ|>�k��>6!ҷ�76�z�����tŕO�s��.�����'n�tZ�=�|b� 	��]=��\͢\d���(������F�C��랢�"ڡ�}��s\=��@����A�	��)tO�c��?�HĮ8�G[3�aװ �ș�b6k!4�����4��u��ۖ����I������P��a�9�f���΄�Xۢȅv�����\����l��.80�;������NDWTv9��1ݾ���$8��a��G}5�cM܎'n�÷[�O�:A�c�#ۈk�i�9{Үm;�D޾���Y��i8)����7��ඥt�TK��L�F��P��?�d;��h5�}�Y�
WRJ��mz���"� O�Es�g)W}c���L/����F5��c#��~��
9��%��h�I��1�F�$��E���(� ��Ħ�&�/ ����v��J`�	׳��3�]�3'%�������{}c--��H;�9�C&K"q��c��ʆ��8d�dt�������	���}��~>Cy[�k.�i�N���=�ԥ=�~�N-�����5F�������8M5}Đh�o�i��{m�,~�mW�Y2~&���L<'2�nY�ug�Ņ�-�������w��BtDck�EWgV�����N���q��#n�u$����M�	�i�$8֘�0`g�|	'�Ԧ�T#�dݴ<�s&�D�ƺo�����IAH�r7�5�5�6�B�Ū݇��n�>V���bw�����L���Hy]���T#��V"V�!}V&(9��I�#�p���}@�]�Ҫ��F�/;v:�� SL����C�E�C�I��X}&F=�L�:Eژ��ӛ���+�w�kB���Ę2�Au�ر�E\;8F6*| <�:'v*�j���
5�l�4�ߢ���#"���8>/=1���F�����8���'q���V?z��a�K���6n�ܱ-Б-�5c�K�m����ma��1������6����պo��b�|/D���ӛ�dUiۤ�����*6�1�8���Y�x�+��U�y�LK�rw���{{Z@�3���k�bv���7ꑳ�����%cT�9�Y�Q8V�AZ��1����<�����z���.b1Z��K�f�A�ًRP����� �z:F����,#������D�Y@ -u[ -�G�G��f��0&	�s�Ĥ)�����N~��][���!�nH0a:H��0�~h��|���&�T-6�1p�%�r������N�+����T��ZN���%��69�"����qޣ3.fk�7���':�i�� �g��9r�y�}�d��|�ќ?�D�#yH%��$��g,uyq�H0�2���Tum�ox,������=.�66UՊ΂�������0S ;�vw�V�c�À�t�}nBź�)�~(���zm�~�ϧÇ�i>���n�X��?�=�DK��=����D�`����n�O���O�s�O��S�� ��qd�n�8娐�]aal6JR�C����8�8.��WLWj����qS<qt.iHȡ%{���� 5������j(�����)�#��R��_w5i@�l�W^'���L޽�,��se��;�Pdi����l�84J��ݟ�n�u���߀�Wd��J���&�����aƵ��IZ�,����lJ��M�8��h���*��ˁm��j�J�m������T�~�wƹzjL� ��v��0}�;?Hw--xDDQ�p���jºJR	�m�.���V��`ˁ1սE�ƌʅ����!��� P��Z�W�M|�}}uZ��ҶA?�����;�L�{J��ô`l��R��ᎪQZ��9�7�\YN��]��z�Kd�7��q�s���n���-A�����t���0!1FEN��V��bYb�����̥���f|�8�,%��?�߀	M_N'S�;��~�@�L���p1@���y1��1�k�u�E֗��7�2���ם���\7L�*�;4�nB{����u���0�� ����`j�"'��lmM���v7���:5����nn��A<2X���p���)2�4'��ؠ�bw�O�7��"���Nt|O�����y���cl	���W'ɀ�$UN�}�xg�{,�I����e{؛����e[#��5�T/o�i���~���mE �nM�0��RNY.l3q�ޟj`�ks6��U�R�D��y����ɚ������;��=Ʋ���� X�f�kc��&����s�6��)��Z��_�q洸�O��Y��tNZ�C�QvTm>1���L4��]�,�c!1W�d����G �8��4�}�h#Î��y�M��L�Tbև°\(%�O9O�f(?W�U	&�$0������y2���a�V�[���iLd�{���y"�a��>����l>��Qu�rB�k)fi�1r��]��m����_��1Z���d맿[�-�o�	��G��9���6o���u��9��u���Qi��6�:�%�p���X��X	��G��l�:)���56��iNm̅�aSpP��&Y�����W��:�me�iTO�O���Dc`�s&��4ZM]��^�M8��,����#���B�Ŕ�U�����h���+;R����b�	�S<����S,*߶�	�b2Cj|���"C�"@�衎!Q����~R���c�� Gl;�,#�ơ�-%X̛��� u�a���A�P≢�Wl�1m��Fk8�kꘖR�h�l�u?��Ꙫ��0���$�'o����sM�T�"�3/K�w-��&�l��Hc��N�<dGG��(���4�c�fz}�#�DƑ�b4{Ź�@|*�tsD��^0�����D�m���U<�ei���:�N7~jT��&�v�l��V�G@d�!v7���V��no�`���մ9h�#�Rj��:+���x��r�������L�u�����H�_��fd��c�w��:����9�W�"��F��v����x���!�X	,���G��s�Q��\����$�(,�������	��E#^[,����y�n�+���{�N�q���	]н0Ѧ���'@����5@�K���Ԍ�򣻝�y6��Ud'���L�4�_�I�6�T�H�GS��ޓ��dAj����Ɍy ���^Lw�Sk�E��u���(-���PG_\�c@5N�y��T�"!�^�R��{9P\27�� �%���Oa@��dRT�T��Yu�Qy|-5T����^/�ncuc����:�~ʙd�T9!y��o 	��M�J��P�G�p�I��י����kg��l;6Y�Y�hc�� 7jc6�@b��N��"��=�(���,3II�:!a�d�6L�Ʃ�6]1�*͗�S@!0�RI	�lJa�C��6#��x���ڶ�vWLmg�"/2(*�`�fo�λ.]s.�+1�NS�I6��	���2,I�1�h?h/�Fɸ���z�a53KW�
w��S ڪ��w6��Dj��Cg�$�ǹ�(N�ͯ↹�X��H ȏb��~�����v��u]J��?�*mb�*&{t��^�$p�VY�`��Z�D�����b������<1��%&��6h�+��v�?-x�*�$�� $��U�G6&�������ƍէbH���3�4?LJ,����nm��q#����z�<���
�����&B"'��D��F-7H��\e
���2[�,4����&��M�I���d�8R������h��_m�ڦ���^6,˄@�͗,�n'�D�*�=��k�����{�`�f�I����7Y�o3�x�v�!&s|G
S��<���B,�?��3d��gu�z�h#�_���:�NZ�׹w���JA@W�����>K�M�%��
LU�ak#[� .����� ��w&^d���=:n#~8FDD�SL�j�蠋�(͙b�e_>��5���I [6��p,��H�3l�d`r="s�Y*dN L�4��Q5�P� �؄��I�	��� ��-�6L:�L�w|'���7\�"N��p4L+���F���~�9'@��.ʄ�D1e�@�M�K��X4nr-T�`_�җza ���}��.�X\1uV���e��JX����[4	ިsҘt<>���Ÿ��Q�:�d
�\ �.TfpV�g�b�d4���"�o��!���Wm�x�0Pi�k�Gg��c�7�=\{z�ؘ��y�s�u���=�s/< �c����a�3�换�:HsUx	?%^H�V�39͢SL�}�*Tx��N��<����Jh��s����ў}$[�Q�E��A����V�v�C!:y�J�W(B!���Nm@a��%���4�Rf�n�*�Z)��i4��J��:9i���������q�ur4=;�A,+���B̈�&#���ﴝ[�ʄe��is��U�?�J�߰c�븬IՕQE?��MI�`*�I �P��1D��K/ubI�a�tyw��D��l�3��n�U���$g��];��Wz�>҃I��Z찡,)����{ 'L��Efx��� .��2/MX�z�!�uW�ut8Z�{Ǟ����]w���;��{�ңO�(T�~;�,�n�u�����Jc��Ļ9���F�cˈŗ2�N�5OS&��6�2��#�i�c�� <�@���vO&��?��k�d���Yp��}əyUO�j�I��[͊��ȅy��h�P���Z��<g͑���y�g�bF���h�����o����J�D/��H)�C��h���Ѱ�.l�wsrVd�J�&�nl��=ת��Z�s�x�Ɠ��̩����9/SN��Uk"th{�u`*�L�2���O�y���[a͋��U�pL̐����Dm�\1��_��w�t���������Z_҆b�r��A�=+��Z�� ^1t�h�`@͹�.�@ c�f�TS�r�0�tSD��9>�E>���M�|�3��=P_m�5Z�|I��7`̀0�O�yL1)�T�0��"���?�gΆaҔ���=��H=y��$i��E����4�>9��(��=lz�!��*wZ��o�!��p=3٢�馆9:[�x�*兺�i�ôL�1��U5%�yO宭~a�gp��r1�ln�Vؽa��k���4*5�M6�Ϯ#^��mA-nsU������_��X ������<�)Ô]8�T#@�TN�p1�-�-^S}	=�y#:��(�I��n��U$f�Ţ3�OF4U�m����ǐ�-�*�2w4n
[���A���u��l�{v$x����Mc������8�Ԧ(%R�b�k�-ΐ�F���A>��Κ���[�>'��aqi0��5�}�vHEgf4G��(��C�x�|T�b�v����e���$�b��4� �8h֊?���PR�PÆa�M�UeF�b�0:α5�t��b���Ƕ���~���'x㼃��E�쓣�ǐ4�i����dw�_��88�q��ȯMHf�O��O��O{K$���o}�mx&�caC>�M��lBm��ZJÜ=t�9��A��p}H)�4 �L���Z��rvR�+��xQϣ&(�C���c4��{�v���fZ����V�@?,�P6�ҍq���߇+[���C�l�~.�B��}u��3���������>�q��w ٰ��qb�E�K��\�8T�W�P�{bќ�؊�@o+O�l�1ck�sN��b�v14��u v�k�|���Mm �JP����t�N�mJ�FR2�χ�r��gK�� ����p�M�����][O%�b>�u_�y��.��i�y��z�F_4)�N*&����8}�C�|h��ƽ�&4X%��)�1��Nt�� b4�|��^�����p�~t\WK#=?٤�7&X0X��7qM�u�>��P��z���1Os��ԛ#tA�ⰝB͑(\<,��y�*Oi�Ǎ�k�j`�H!l��^{�Ԇ, M2��t�M�]�~x�9������l;}�:JٹAhW�υػ�4�:����g>5��{G�G�Ɣ���{�d�pZ�i���M@�Q{Y�\�,|�(h�-��>s�b`@oB��!7�`�@-�i��ձ�w��;M�[�2�����0}�4�Ʈ��Թ��&�'`�)�h�ąцmdJ�7�i�;�e�.�5=�6�!j��LE��:�1BE�]�o/�dX<�;�V�X��~���u-mm��[�&p�K폩�*D�cE�m��+�q����?��7��j���E�:��8�4�ά��-�e�6F�`~�F��ɨ㭳&�OxM�Í�!��J�]T�L}e'������\rI��)4�̚��[Qsh�6�����g�"Lt�A�mW�;���zo��]s��*�$����7�ɳQv&Z4ׇ)��DS���ֱ�U)�s�q�O%���\7?u}�R�� <��~2�Z���:�m�V�7~��n�X0�{eI��#�M�D %)�lXn
�D-X&]]
����w�ˁV=Q#x0������XY�9��`?���A�Bw2ؠz\|�%�=g�Vb`���8�(�R�6�Z�,�(|�0?�[��f���+uw��g_l����R���{�t]=����h���͹�ۻq��c9u�=?-����Ѐ����f�O�A�T6��}C��{��k!=ɀڱ֣*RZڶ-]x��q�\<5GD�AJ���j�ʆ�EK�L,p��DV�A,3o��*'�5�x���4�bW}Ւ����2���lLE���)�)�9�Z[јp:M�a^����0�8x8��ƺn�ޝvM��R�J��봲dp��!���j��!�y�!��`�~O|�h9USv�����bP�<7��s[�;}/o߾��J��P��CM �φ=�e���w<CRp���ɚ� �u�z�f�Bz<D: ���������V�4�V��4�;�U�
J�z.:c7v��b+u����\�zt���+��Jm@= �/�ls���NX�ֆgp\�6R�̓��IT,#���>,���<�y@[�^�p��|�/-m706)l��ǾKҒTɲv@��L�(;�_�C<�t[&�!5aOEV7�\%�fٔ�d3Un��̮I��,L��t�������Ҏ��Vnj ���������Â�ۢ<�p�2F�X�=����x�׆�g_�3�k�N[-�_Ӊ/�_a��h<��zի������b��y	��M����Ǝ���Ƹ���Pg-q<�1�VD��Ą�cFN�R���ņqİ�c#�����H@�{�1���Z��G>��gs}#�B�S���0��t�B����4�)��ͼ�YX`���d��VǦA��)�dߙ�����wsY�����&��h�Mh�^g*���2�u��D��J��##b4J�d���W�WݎKQ|��F�_��z/��)Z6m������1fz�&�+�w;R���=�*�T���(�6����i �Q�����������t"7�»g�]�*[1�JЈ�|���&��;y��E�Z4f����/��/��U�w��Ƅ�������Ռ��,:�x��Ԅ����,7�gΑt���"�D�v�q�^�d�n"�5^��].�=u�Q�%z�SVY�,M&j^�E� ]4@g�k��t���Rw����NZ$��>O�:�l#;����a��`�k%{��D����dV�K�7�ܤeD#�Q�����%&u;Y!F>�ϭ��ܡ�c$�W��@�k�@�=8f��d���	��O#�@��Z��f�H��/��<�ǔ�̟}so�L��\J��d�x�4�Uڜ�:�����»/ w����S�{� �N�O�7\�%��漺c	ӹ��8��8����@�<�W����^���?�A�|���p
 g)�J �u��i�J�H��	��c��M�O�9"�BMg1��`��6��K</�=n�Ȣ�jL,�E����t^}��n7��G?�̤��o�V��?�c�H&Z^q��F�͖6=���m(*�Ԩx9�l����u9�B�<C�3����^쎿�|�QAP|��i����g����,?t���qӪi�X�r��QZ�.�=,�Н��۲�86�3�̞�&4������o9K�Öp�=*\P�|�|%�E:̋z���Q���'A�.�.��-��R��[�/�4�yf�h���%tt_ڴ�L�:�K�����I�'w8I�X�g7�����L�Ns�\�C�x�.,j~ǃړ��o�Zݸ���x��,}��ż +��a�~����{i�<G�V�g�o���-F��GX���7�A�LII�-;'t�Gi�9�	kZq�ZZ,9 ��Yeɟ���1�ͅS�6Bm\&P^c��̚�����o~�g�D'���
��^���ڧ,A�h�K]z��=�n�s�$%�Λ(;U&I��p��w�kE�Ջ��zS��'^���v!��n���t�Ъ�g��Toq�$�&�y��=���-��>��1Eԓ���H���~�k���yc��s��`S���v��
��9ڀ�F�^�"�g9/�}���ϫ�ql
ӈ�&��)}?ޫ�RM;?�Fvg�����L$��g�M�lM�����{W���4(�Q�m���A�Q&lQi���%��}ዼ�e� �o�,�ʠ"����4qq��1&Ј!�Mws����C��uߟ]ߺήڻ�34���tU�}���~��o�L�͂�e���%�}w�Y�l���#�_�ş�m=?� ����;�JzH:nS^�G��f��m���꺧e��X@��>T�	��I}j=��'�i�K� F�*�[K�1.�H�"`�#�=�;-��Ս�S� �7/��J9�tL�]�=���:���j��h���§�?��W}�W����� �l���=Z�a-�*b�����P��А�I9o�sp�3$C���%v�9
6j���YHK�cx�+W�){�=��ǚw���}�io�:d��VN1a�ӈ?����5f1-J� ��u}�����8�1�ڎ\�1tP�k���ph�f���h߻`r< ����1����ZF�����@�7�ɧ���y��9�G�gl-{+4q��x�w���K�?�5l#)	��d���7�Q_����m~�����?�áF� �����-�j�Z�	�3��w�l
�E1�Fx~�NjEc*�S-�������,�������(�n�A�,�n�<�ƪC������,�^���?��r�1�1�a���@��k0�<c<�}A0�LdDk"c��D�0��5�yM�,Lt�-��|�:9��ps���
/ԍ{���%�s\ �L���߫s1�k�ZM��v�=���:4�|��=~m�	>�ȣ}Vނ��*am�o�$(����� ]��DR@ee�עд��L���M��s->��S��a�Vh߸�bΥ�+�@�i�V�㈾w��L&�X��|&�'�-:����8z�� k�ױ��(���h�=Jm�[�='������c��1]ڥ�}%������������gǏ�e���0�X�H��������{��җ�z׻�W��U��^����BQ��:��g:o���q�d$�ϩf�!��x.��|��h<����Ɂ�s� �O&7�a�j���y��"i�9}�>�:4a&:x��v�=��=%���:xC��?���q�1ji��'e<�$��j���>��p��Ӳ�r;l�9��F�h?�X�z��Ds�-?WP���1Y��QےSЄ�x�䕽�g���|ڧ/O�>;oww�L�@Ts��#uw<�Q8�_�K�z�C���!L���.��km���\�7kx$Ր���i���uԴV�D25�!�$�M(��Arۚ�j��&9�右ԧ��&��Y=����ܝ%�G�8Q4Kj��К�h�Mb	UcK���I��Ej�q���ӂ�j�7^?S���}
D� �l�%�@t�l��؏�N;���4��x��;�A��a�CA
l:�Zt 7@ȿ����1�wc���xy��έ�,+?QeNy:W�T��A����tB~��4#t��9�����P L:~��++�k�d��%l��󶯐F=��bҁl7q;�q�N��ϊ�eT��+�Ep��{�찱h{��h(�Px{�U��bqXwb~Ѓ<�=�Bq��;��Z��p�l�V��ս�����xf�+����o�����u2�E�䲬e򢂗א����w�m�L��woHmE���JE$�;񼎜5���j��<���g֒�s���¡W^��J��h�v�ԕ�;�I*�}��M�����1�<w69���4ۏ����;/}�{1�q�!�`�h/�%�W��v��3t��*<�5nҿ`�t�%T	 0A,���J��i��dMx��Tc;+� �^F�X|�+^Z �����b��H��9��z�iDB=hh�uZ�	!��M�T8a7_t���/���MozS�����z����LQ��jٞ�w^=婟��M�>O~��.���uZ�b�M�	�ޏ�&͕�I�����.�&<޽��~0j�ߠ@_�}���{�Gy��j�m8]�:���e �յ� �~}/�����ﷇ%���b*�e*m��LV�{�}�V�Ϭe�����;�ɽ�N����'}��<n������9�M�-"���֠u/4�3�o����MGM}LD�g�g���~پe�|���򓰧r���w�^	��G.<�>f��$�>j�_��=Kz/�˒����0w�F }��8yv��P�x���ȏ�HyBW��ۿ�` �,kS���Ll8�+�`]�h�j����x�Mr��K1}����i�l��F�0Ԉ��-@�p�7m>��Z��08՜h :�����9�A�\(4��_X.╯|e�v��_����Mf��|�ה8a�w�աL�t�!�Xj�P���o/IT�"�c���"���m����H����E��P���nF��{:��4�+�t��Wڍ{Q�`^���)4���1ͥ���̛e�qn��/[��2Z�N�^��j_d/~��/9m�� HH�0�8��YZ��I�i�b�2��h!3�.�k���~˷|KI�b�������_����q���Z�8H0#����#iK5^1�s��(�;ڊks'�:���S1h/<:�4��0�c6�/� �0�y_�З �f��	W���X���r�(/��hDk ���[�Z8 �6�5X�h ��6���P4�-����/�i�&&G8/N%TƗ6���(lo�y��h;�Q��+���ލY��P�	J�ٞ;�5�5����.٨�[����KS��C�:�/��m~����e;�Ns�C�oM#��VǶ��9�~��eJM�b;-@���D�Mjg���?�Lk��U����#:ɚ�ʦt�?������</Z1|1QS�IF�Xl�yL�.�n�������n�c���h���~���Hџ�n'eXSDK��~o�-��xz�9�yn����U@5�Qn�tP�����AepM�BY�$�O�tb%b�"&��m(�#@�Fռ���a֧E\�(�X�Nh�=G�$��L�}�Jj�Bo�8�+�X�o/i�MS2�F@_�z_�1&K��q��@g5,%��k��6j���tr&��[ṿ��9���~n�:�l���f���f��c���|�*R�s���T�N��:�Rt�3��"qȓ���F�3?�3P���"w�A��:d���2��5f�N��҅k��v"<ҡ�mw��s�E���������~��>�O%��s��9�QXa0G [�4n�B^����ĺA��q6�f�GkF[��a��m���Ȟ�zm���J�-��1��b����%;���(�4����h�.�6�������<���L����G�5ړ&�0Q۾OF��IC�)��t�3�U[�di� �����'�(J���SN��c\>�
Se�c3U=��{�iE��v)/���X�k��et�d�&< #��%��ǝI������'A��zqqʸ��X|뫨����v����%�΃a
�����8P��z��Zx`V!~Ҙ��h��2��f<� �f�3L��c���Vɧ���������a:��߸D?L�^�-�/��{p�H�f<�U���z�Rf���Jv�25rѧ1�b'[)������Ak�{�5C�E/�C�r���]0�H)�v Ϊ���d6��A�+�*C���=L����0�Z6Q��M��K��,������OxN�b@�H�YZ��BQ���8���F�P�_��Хh�p��x$Z�֋�#JC���fm���a��br��,$�y(��)��B�~���8��|�s�j���%����3�+�n���9�`8�㏼[֝��u��M�މ
)��P����Ė�:g}�>�3���[�Þq�E30l pI�q�ŰS�
����WO϶��%p�=]X�e���	_�����r+���Y#�qյ������I**���T��SW[q�G�s�	̂ߑ���6�Ęm~�������6܏W��CJ��35�<��qԁY`ֹ�9m`Gٔo���C�?�UN����S�=�Gn�r�͵�5�>�f���2n@$�U�m�����0����
���Y�*��*H��Kj���gL�I���Jl!�����"��+�q��Җl4����Í�q6lٛ��sQ6U,!-�i�ϕKI�a)�c�5��4SգNЧ�r���;��>{Ϻ�p��!eF=���xnk�x�*ǷU��T��y�kA����P\�7>��ris�NI�	E�@;�O���	 ��9��g֥���!:��5�����3�#�d�C�ס�}`�:�Ǉ�qR+u�T���d�)rKj�5a.@g���l��$鷋�,'ʃ�ڎx����)1F?��	���5{V"ߢY2��t�O;-{�!fK(��]a�rl��#�mn�܉�o�yE����cW�����)��sM',�4ڥr��γ�x�JTt�o�(��Ӷ=ǳH�Ů�N^��]^:��c�T��������q��,0�K�?��w̝Sr�����>I��G�N<��?h�y+��ޠ�V�w+�![�崒���~�ߗ-���4��΢m6�|: �z�W�M+<����V����!u�S�~����I
�I�$��5g�4��ٖ���rF	̫�n���~�����RGc(�FU��~��wV�
M�,@|r����b#�$ d~.�m�(���滕�|��y�vS��*�=��׶�x�ss���5�+	���^u����oAz+[yb�y��e�����d�9�xf^8#�ڱ�f�me+[�����8+�x֬R7Q/R��i7�};�3k�.�q���)�-'���<qe�OhU�^�y���*���	�N���n)H1ۛ���>{��|�Q!q�f�el^Vg2hN��5Ӕ���6_�Xd�#��B��4P���m�t[9��s|���*ӯ�`�
�O9)�,���DZ�s���\r��N�:���C$�`��kȝFΛ�h�� �i��I0�9��w�sS�3� 3��td��c�M�����='\J<��O��Mg����+[���zG1���������9��[X�
jf�X@�x�6�ŧ�\�L��CLY��j9S\�	�)'i%�����}c�yN�e�b{�k�Tw��϶V�v�=�ռ2=xUM�z�;	\3�vG#Y��y���!�o��3=9ے���Z�s/::��r����ֿ1}��`�G��Ӿ�uuz�v�;Z�԰�O�[Y�F��Ew�����+��Ȁ��C�bn��dCԓ��6<�n���f�]F_�
���� |�y�8�:���R�:�cV�����LA��%�]�o�9ۮ��vzזF��*P>�O�`O3vΫIg�Zֵ3����cb�J ���Z�f蚒L:��ӁUVU�������pV���R�٨�����bSv�����G�8_W��Q`��Ǽ8`�N�!_���`�bd�d�[�˕�MZ��t�ֳ��|�C*�������x��ǣ�2)kJ�,�L9	���]{�8�D�ʸr��IB�����.I�X��8z'���ˤiR����u�[��B��Y��ZH���w05]��������(u#����N�v
��W�."�[*3ۚ����|:m�����H���~g�8ǻe��g?��e�^��GTw&
�%.)�p��=��x�41�G�����5A�/��//�Q9�FB԰���J/�&���i��d�{M7�,̀��Ȫ���4A}N~2���� �-s�%�U�A`�
��֝+�iL�֌�ɂBtn�$����Os�ӊ��|/bXn>�q�VV������g�
l�6�#���T��d&xC�]�Q��1�����e8�vvڡ:P�}4�\L�|v���^���y����BV%�C�MHV6��8jx��g�8��]3���W}U���5��k_�ڢU��~o���		`#TB�o�x�UZh=iO#5�X�l^7�s���6Wq��-w��=��K��w�d?���bCaj�J��~�p.B�c�t�*Mv��c>�Rp�0U�jk�*��Ɗ��������+|��e��?��?-@��(s�-Q��������F��=�tI�mt� ��؎x6���lY������K��-���4��<�J���'�̆}��^_Zg���AL�p}@͘	)���v�s<��NnX����ҳR�9�4�yMM��4�$�z^:��kgIĴ�r���E0�m2��ww�I�Y�d����}�Y7�Wi�g�\��������h��'4�t�%��ri�_6��P��$:��������= �`}s}�oJ��:}Ԧi.A��Jw�	�N�CǰR����̧����R�݊���N�Gx94TL^��/yg7
u ������-��_�x�7U�9���lYM#
�4$�cʥu���x��G�e�H~�����owQ�3��e��ŹG���zCG�Pw����7�U���w����y�i�o�9_;p�x�\���_�=��X��F�<Q����;w���j�75Ԛ�Y5�7q��ǿ�����:Kd�Eܟ��`Q� N4Y6����_��%�HG����Х/y�K��P����(vL>�x�q�A��<�X�+��+E�ĺ�6�:B)��s�^��3>�h�t�������_~xٱ5#��/�Ơ4 Z1+��ԅQ���c?�cE�������5�{<q,�����tXzVW˨�ض~���ge�N6�/v�M7GlY��Lg��рp���-F]�-��>�V�)\^S�zQ6���iL���x���	��l�Xn�Yvʘ \��&`s�L�Fv�6�^�ٕ��b���^�κw=�w��)�=Yx�S��;C��E
�!���G������@�����.)8:X\��?s˘�l�c��������n�)~�J.()�$�%�[K_���
YJV%��5��?�3N_��]m�F��>�s��������׽��2�%�k�7ύs�x�[�R��s"`;%���/,�g�b ���MHݐ�cxfϷP<�>�_��]��3�\��~Y��\h/l��áŲ
 �L4M*�&C9�2��5�8��b�¯Q�cJ�-G�dr}���+t�7}�7�p�n� ��|���>�w��Ґ��W���/;-�^5;��y7��zf���x/'��k�:��4�vV��Ѽ�9[܏5�3-G�_]�X���w�����~��q�i�������4%���]:&�Bq��N��?[.<�fm�N���:ۦ��6�� yw^0i�]m������,���e���a�q������������rZ: )!��DY�?���B�o��ļ���6E����j�*HI
RF%����J:�yf3}���v'�|n2̎���:Z���Ԏ�Fay=#r�C��ъѦ�+�jX���.8N��\�F���<��4�м���备?��惥G�4�<
/�>N��4.Z1�n��G�����ſ�e C�9\�E�x��ye�i�@��݃י���ʻ;�d0�H�{������®C
p��8��i�N#�ǃ���Ԇ���>���]���+�9$â�@��]>��� �N[���f��כ��N���V�!C����u�$w8N� Iڒ����zf,��Ay5n5����C���h�Z��|9�w�n��N���]��M~ү�- @�~B����]m��=5������:��J8�981g9�t�����__@���/��|M�������=yN�%�{��9p���X&�:F3��4�
$44(N:�o�UЇ�@�pV�*؁�����}ۣ�f��~gRUx���ܣ*�s�Hh��X=��̎1\�kp]V#���X�8����1���t��_G��L�N�m��k
p�A�l� �u���ɴy���Y����On��>�\��)��J:�n4���f�j7h�,�\2ل�/FJۃ��M���#�8��a��Y�ni�䈻����W��z������>�i��d�e���Q;�l�KS���a�8q���1��d2��kq}���o~s1ɐ�]l�@r�����jS9/X��"�����T�k5U�Ѽ��C&@e�WF� �=�P���8)#��r���� ����/��������.�>	@73��*����:�ZY����H�r/>�	^l����k�q~�tD{p�i��Og�x0CC�/������;�Q��2H���n�t�����1��A�P��4���e8��t�<�q�7���{�o���sԻ��2{��g~O����o?e�\ߟ�ĕѸ{����f|�����|�k˅����\�
�:�����y8f6�μt굝	����{�m���zj��]��|b7Jz���μ���Kʹ�׉Tm�֜焳�4����O�����51�c�#�a0�%���ó�w�$}PG�lz�����ڣs�߇
�o�D5��\t�Ч(C��I"R�ab���y<������*��+^�l�5쳨ȩ4�ǻ�#r^h�!�ͻo���B�uhC���]��`ؓ������9�;�Q�K���R3���0$)�U5	����1܄I���te��il&4�<&/��{L��FE�̣%��	Z`�v���9�yN�_���=�����z3z�Ϛ��?Ҍ��E���pʝ�v����f�x������
���9��X��ۚ���m�#�q���'\9����֠8=:�|��<���7~����4���;��4�?��?o��)f%m�IY:w�(�3j:Vs#VM����F�߹�2�є�������KG��[%O$�w���]k-��P0���
���j&5���� �;ᤖ�xp14�
�bFF�E��TԸ4�O��O���~&�@�@�p���Nk�q(�߶�J���f������E;���bAx4���X�i�H]t���<��Qr�#�K�A�5	��������w���~�����?����K�S*��iY'�����9ٽ����a�했("��rOs���6�Gn�kݽ;P�>�5�����DUtϰ�<@�eA <��jċA��y	q[ x 7j������aG��l��~�fr��4�w�^�R�_���i͍eȽ�������Ȣf�+>����t�jN�vP�Ŕ�İEǄ|�� ��2՟���Q󹧑�4��,�e�8F�4�Ȑ6R���<4f�B���!�.s�����G ����/�Ғc���1>0V����x�:qG�v<�� 	��ul6b� )�����ީCv�"�l�ߘ  ~ʻ�1���^}7�19'AY`�U�@t�\��d�!�|��w,S��\jr3��t���u2��Y�o�3��/�� 1�~���^������ ݶOp��xgtown�M8*�o7�G�zFɹ�l �f;*�C���#����>�eQ����B��17�g%�n�so�'�EHl7��t��$����7�a餱�\��\fB��aB�w<�a3�ԈV�9�<��"��1�E��v7X:!���Z�GbÛ���%ݘ�ٱ.06���s�S�����^FE1f�d�b)�S
��/@C���q�w͒��J�»�1,0\K�� ~1�LfW�y��� 'k����d�3o��t��:�lR��S�0'���,1�K%�a#����?��������z����^wa�&�>�w��J�/��Bw��x�1��]�7ˊT��g���g�����w�%��j^��� ��r/�'
1�=�)�c\�3F��YF%ԭ�u�6m�{���[!�#�5^:2U9��s%�ΏԞ3�že ¶sj`ϛ2�uKԚ`>_~��+�4<FM/#C|��}k��e��mb"�����$ţ�{ؖiu�����?#e��/���:���A4M�gU�}��h����3�5h������0�B!��+�����@�ö3x�;�b��h��ۖb�c���}�� x����m��ѓ.<Dmr�8�;X��$n�JD�X�G͠�l��>��lP^NS�I׃�Q��`p_��t�f��zp��C4K ��d-�bH�P�1�GC�D[�[��-l.\-q��$`bu�
�nw1-�=��Ym��g[��ܩ@k�Q�f��iw���s��<���!�u1x��>����Ӄ��6?�aT��}n�V*����i�_��q�#�E���J�vҪ��g�#Z�z��D�tg�*��E��`	��o����A{BG��K��E*p����g|�gM8�\�
k���f��Nx�N�����r]�cn<A�;L����ދ�[̎�����w}������9 �%-�����< �/%���h��?���+_�ʢ��Rq-@��~��=Scs�_k�7=1j+�K�r���d��~���Ƕ2�Ƌ���
��
`��j��<˵����h�]sZ4�/S��� �{���(��gy�����֦2ʡ�`yέ�'����9c�gE) ԰���ӌ�Ur+�?�Ll���m>Ǚ��l2l*��N�U��E��!dFڀ�mԎ���}3]�������Ԍ2�j�M*�:8j��j��1��.)��������F�x&�{��dg������ާ�|��|�ou��e
1�B�X�,i�j~��p�,��j���� M� �C?�C%<��D
3�S���?��'&+�I.����h5��w��.�5��:Zby��?�Utџ�����= ����pˍo���FK���g�9�3�-����V���)�j�L��0I�0.+��>�����2Y�{�[f*I� �IOhp�s3��J��#�����7��lG�-?����׼�5K��Tz���$�E>���b�
m��m��K��xi�Y���+~r="��{ǳ.(tp�4���`��J�7�s�< �����JQ�?���^^Ƽr�L�/����g�'�Ά�g��w<�@�Ώ���7�����*����'xȐ�*���w��;���4���}t�'W,O�TKr܈$��YIY��~�k�,i�vI9\�p�����V�yQ�0�?�5�^ĤP$8�F�q�d��i*譺f�}�l�xUƁ�pnJXg�7&ΝP�Ƕu�:�y'	tL���	��.�i��iZ�e�#ڌE���T�Q;�ְ�KL��{<�[) ��Ǳҡ*����^F���3��+��F�ʚe��D�v�],/�;�|6o{p$	bV�B�������i�����?�3������0�LWE g'?\ +�8mM�7�́�F��1:�t��y���=�I��a�mh�ĴP��輈�y�c���%h���+�2_�K�`1���G��iz�F^*��c_��p��w=o��%�2g{�U��YD��@ƕcV�ؕ�BVQ(�~�v�"�P;M�0��a��t��r����n�\f;�FX9?�#?��Ji)��:pI2L�V	�i��*��H��b�p�n@��P���Ң�br��Rk5ᲂ�g���U��'�������_�P���P�`i9�\�T^���2��5Ip'�k1>��P{p��1=���P���0��h���6�`�4�u��VJ`t�`;4�v��zƢ��h{��}�"F٠�>zTz3���db��n�i�7�V�!�b�!�����k�.�L�̶\�ӆN���r�]@�	�x31�	Ř�B2�`���w9���y����`&�P@m �$�[�p�EN���#���a�o��9���7\.r\��W�W˸�^
T�b����厵��� l��.#��;�]�c��e��y�}�����>�++�����e/{�T*��@+f�#�5	-�jD4*�5M��#�w������YrţXƲ!���@j�\S����'��m��?��&R�?��m9���<�v(WIŴ�a�ʦ]�UTø���7:R؇�rM��x`GM���M�0T�,��5�=���Ti��J{���&0ƨ+�1� �L@��z�s�*mRJD�L��ա���=���y�UϙV���z��h�EΒ���������^�e,o0j���Z�]�\kP��0���;w}�8��Y~�t��MтKxǨo�v�.+&B!Z.��I%�C��$�����,�+\H4�����E����y�M��AZ���k��f�[��҇�;)tA���i-��I���P����n 1�;]��d�,
1Q�<�9�z�C��@It`M4J���I�i�w�.f;��Ш5a�n�!:�se\i�}e�{��P����Y�6��&xL:�,���P�K>O�}���j�h�W��ssFDʂ�c��]ES\6�՚�����3ӄ��p���3���W��ʈ��s2c�3Q��Q{GjJ���Y��*|��M����琚�����UERyO�,������W�m@�O4_�MF�a�؋�D�Mmap�Z@֬~:I�^s���r׃�����Lh<9 ���@,�cxʺ�آq.�!6���>a���b�y�ա�X��N�^�>Ԫ�k��$�/�|�ŐI7/��6r�Ӿ�p�G[�|T�cvx�2�}�G�N�p��ֆ}������ߝ&m����;A;�]���7�H��5��^�]Ԑ�� 컬Ɩ ��S��[)����T) `�A)(O���ݖ9��Ox��ؾm��Eu��;��5�ub��2���;F��
E��ǭd��4G�z4�A�6v���vz�����]c��!"�-������_������DD�������DN��vI��(���J9���c�t�[-z��i��@� �7�םE�b���,i(5d;_��E�>L��:�Nt}
P�������n�?�9}bF��`::-ƣ��8�BS�`��{��y��OV����5̪y{-�L��_�М��:7�`x��]����&�f�qK6��k9p\�LS���˘�����s�H����0�����8w�ü�>�m�'_,�Ej�#�k��r�X����/[zxe4d۝Oh_i�:6�󜩮NNk	g(�f���]���4|Q-"'�I��z���8�?]�y��U�g���}e���6��� �S>��T�ѡej4
c�N	������ͱ�bg��eb���ye=�G��e��KIj�Y��Q�����V���gu(c.5r�F|9�etD�\��2�@O�i3�ޖ���%O��h��q��C��@Q4͐�Ԇ��o4oz�p^��#��Ϛ���y�� ���i�4��K��K�c5wK��S�`�������\��2�����bD�h��|&�F�  ����ʙv�K�#�A�I5O���%��s;~�0�q
�X3ƒ�ZL����bG��[�8VoV�<��c�;q(�����G�;��lMO{�\Zne�|ѓ<מ��6"W��I�ϲ�O��
7.�b���b��ˣ�~�i��Ѱ��臅9n�,5�a�m�.� \��aw�r���e��K9��n�䖘�8w�-)��I�֤SՍi[+ֹ����\��px��"��H� �n%�'��Lx�O+[ >*�Y��{���;� �Q�[��i����� d?�ղAT�tzѧZ�n��δ[!��!7"M��,؃�1���5�1��\k$�&b>hz�=n]�M6P6��D�"�^�,<}�dE�-o�Š�6�C���D%Tl�GD�FC��v	�}a���ۅm3�I'̇�����/'��B����$B�\��E�d}zɉd�~q�p���=�p�kE^��o��>���br͛>��p���b;�|2� 6����@�����������PD��!�v�����-�(��89�R���;u �R�����ùA��C��b'�\���4�hy'{�2jkz?3�z�j�E�[T�#��Eq�M�}�F�ѣ��0���Y�}�B�y�_Fß��S�-���:= ��5`�~���.�ğ]���xt�˄:ᤗ�#��0~�>����E�r�3���$9ae�o.�KI����n`�������Ҍ���Ck9�"�5zo�Ծ �D�Q	�BU���tgֵqLn��l���b�"�f�+�#��!�����q���06�Ś$r�ir���p���^ic�ϫ�,��y���5�d�<i�����}P
�+�޴_P�r����;ݻ�'���-�佾p�Z��� 0���$�� ��|?n�3 ��T�m�v�9�>�P}gҗ�$�����C�4�A�b�E� &���N��?G����wfJ�����H���=�f�<~����3�K��>w���,��E� ��O���L:�c����\�f�p�s�#<�� ba��n7�`cD����y�~�ﵵ[w9i��]>���Z�����T�<��r|��i!��>��n�	��^�e�|���yNrKZ�A���dY��6\�Or��4f�
�6bC��i/��ݝQ��b��w�"���?���w�u����'�3k^��Oo����ь�ԁ���p�0�@������=�KʳsQ6l�qGjMFG̗��)Q�W������/��Z�?|w��������,?������I��䈗V:F3�z2�u�s§s�<��wy��Z�~!��	��K��i{��/�}�jR�s7'�׺�%�!�Y�s�c	8�6|�½���IVpN���g_�&w�?�2+��"��$%j-T�uP)i8-��VM%N�M
"���m���ȉ <ߝ��	�1�o�C�Iz_Xo��v��m�Iǭ��Q�� ��: �
#y�cް��n4��N�8�s�\{��������']m���4�Ϛ��^�	�V�\����i���v��� O�uϸ�(�1!o	��.�Z�?$34��QҔ��4�����f1n�=6o����������h~Os��f�kÇo,9��l��� �@�X��Vk	�Y$E�:'�13��u�F���@.ԙݥFc���,j�	�j�����#�}e;Y�H:0����ZD�]�<�@&���t��/J�┅Z�BI�vͬ��\H|9Fe�s�1}&u�d�Ny��o���8!`6#'w4�!�)�|n��q������C0o4و	���`^���5���;�+��i�;�=�u <jw�G��7����o����G3��x�B�̺�8�+�;�3��<�#��֯Q�yo�1�='<ҟKi��W���qs}�j���,?�9���^�����Y?!M��:����	~5P����?3lP�H�tq�>Qs��djvu��<��J�El�s'H:�k�C���j�ׅlՂ��B���Ͽl˚]v�Q�~�����ĢTH�����\��K��9?Wj�w�B��4rr)˝���˻��VM�H��M �)���~q��d2e������}�}����
�ģ^����op��Bmt`�N̄�=>lf�Ǔ��mv�����G�R+�x1���f���
��;K�[,�s�{�f�=;��w�i����'�&��u��i�Bi��Y������8ps��䲉�����f� ��[J��Y���L�o|�hC��vI߇��{�+MZ�	5/�B�8 "��\�l�Զ��_��"Y�~��h��
㣎�Jg3�vG��K��M��']QYb��E�1�]�m�сK�7����M�aP���o����(�8�(��!	��,6y�^�]��i�;AH�k#S����D5L�;E��ܝ�N�j~v�Z�쀁Jڤ��N��G�C��I�7��l�[hD���yoëa^�O�JUƄ���3�#�ݻ�v�ּ[�g���M:�e��B�Lk0犝INZE
iS�\���F�Ms�|�n��H�I�$i 5�z�y-a?�HB��%��\���+;�����.�%�8�|������9fy��M�q�9�.�i���RY�]��x_����N�����H*��?Z�Z�\�S��R舝����qK��x�����g>�����MG� ��>��>�������	���Ex�z��M��'�w�]5����گ����4�ɚp�{s;'S��` D�:��o�S���v]с!pg�u�2��R�� x��h�B;�Hs���=�Kl_�lT���;*�w���I�N�E����vJ!z��I� s2���}վV��&�hN��$Qp��U�e���,���_u����[m�;��&X�;��L3������,�z7��zK:�8���g�{g�*��R�|�צ���5��`{�Qv����tW�a��S`?���
ճ�/���M�E{r 2�a}��=�䗣�R��偭t�dc0�͢!�E5/F�d@���|��k�v�-��}ٗ5�����R��S>�S������y�4���I�pߑ�i��'�)`6kv�t����$:���������6����N3ݙ���ʼb�K�q�媜7m{_簟sS�B�m�
�/F%�uP�.��,�:��R�S���2���a����i5��&D��I-+��UϷ�=]Xұ�.���;%A�62�$�$���~�Gf昚r}Q�I��#>na8�����pQ�8����He����X��۫�i����2�aB�)�d�L�y>nK����fo:��N;\4����m^���u ���D@��Q��t�uP�	UbB+6p�m�8��������������rr��. �M�m���B�,��Yq��Wq���i�;m�A7�4�����.���%��D�ᜦ�{�-���=M�h�(�[�7���^���34��B�L���g���M�U��i��U��8`O0������o}�Ȫw�%��:�v��V����,���*Kc���m׋��'}?��Ԁ��s�����)��җ����H��,T�wql��
�DBsF�d�$wJ�e��%DGt��|>k�by���^3� Z(+����̔!�A�3�*������AU��N��1Qu��hK/1�x��P���_~SQo���Tۏ��ਜ�j����̫�O�����Ng�����o~�E{���[��:��;P������������%�4U�<`	8���;8������B�4I*ƶ'u�Be����hĀ1��IB�B	g]xNք��j��3�ǣ^�EM�Q��}������=
Ʈ0�4B��3xd�EB�&�AS)�J�~��_] �M���Ƨ1�\f�1u���[��ǻH=AIRnոv�/���7��^���BD��C��98� p��Z�d�ִ�����hJ?�B*��	㬫�
�ˠ#��a��rŸq�F���o��  �8IDAT<�Tf"ځm���0��[���#�#<�+�u�t�����7���s@@������r�g}�g-CI|�4�.#Tf+[�ʭ*��|�(k�����1��~�`8b(���~"�=h8l`�N��p��ɗ�;:s,������I�LZ���7t2j�%=�{�:x �z�]@j;s��Y��Pb��N6VW>��>8����#/~�~��m8�ʩI������l�NK ��(���r��}�k�e���5�w�,�T�����"�YsM}N��3�;P�4_��k ��U�$�����9��\x�p;u�(���7��~�}�'�:�������Yіm(x^�u�4@�W Z�i^�"����%������s�G�u��	��2ƶ������܇�D��bf�z6 _АZ��V
x�N˄��`����%�ŀ�5˥22�c�j ���,
���K��&��ɧ���-/��ݴ�_�E��G�kK\kF+���Z'"y�	�ѐ��Фx��^V��[���Y�X�X����7��7�r��l��9�7���w|�w���/� �@x���%��_���Zǉ-�&�
�%X�ߌ��c��L�87&6�
�������	��S�_�҈W:�,9�ڝ\)���X����I�z�Ь.�+�aŒ�5��h	V+ N��<��f��ߒ�6���[��V�N1�
�{��{
�����/�b�-�jf�~z�DVN3٪�H�6g,�a��>�]{-��gC^f<N�����S��;���N�"܃���馂�1�j�� �4�2�����_����T���%���|��}]��w��$f�[Cs��L-�bH���L��<uH���V�陕����.q�Dc����J��������YW[�P�Lٖ"UcN�0����:8Y�,���>���1[�m'��A�ӄg��br6k��%���],_\�4r��Y�%�=�43���2���46ǲ*q/�l�]����5��R�[�V/�R��W������r�ŰS��o��o]�����I?��?\xa�1�ŐUƳU�bUVf��U0ӿ�gfg���h|�i���|ҩ���4�~�o6_`��?�c�E����T_�H�p��2كP�Cd5����IK�	w�&�U�LIEn��[H���*c*�"wB�me+`���"�o��-�up�8 ��1�82��v-A,q��\�Y�ĲL'g�s��6��������.�H?��фǋ�f��7tܙF�~bfn��d����0�Y��!���;���<�aú�}jv���G�c�
	�:u�2����h8Hub�m�D)����W =�������:�M���`��q ̼c��=��J��
^bG�p�ω�H���ѩ�d>8(qo�A�b�2�#�������.'1 JL���^J_*�T$�1/ $�wӎ�C�')�/zыJb�;�����A��?��%�.k#wJ�F�$y�e��4���
���uի�l�N7�k���ې2/�~��?�ap�}�H9F�Cy��%b�,�Ԁ�^�{qOl��<�E�҇T���9u� <�L
'Oˍy����J�i���������v��� ��FLа� jf�$8Ǒ����庿�+�R���ჸ�O��O���[��vq�����z#�=k�[�\�$%�8��.h�#j�y�o�v�c,`,���H����g^���{�W��������*��C�y��=x�&�3�����Ek£�ɂ�����;�� �GԼ�%/*�����Z�&i$�<��/G�9߬:���9נ���C?�C�Ꮉ> N�Q�Z:��ِ�ŝ!��N���mk.[꺳��1�u���lǭl�v�������5b�`�%m֬�e����峟���(ו�����k<C���!^��6��]<'\d�� z��~�l"�����R��*`4/'��Cb����2��|�;���w��h�hŖ�C�u���3�3���@�u>5��'��� �I��饈N���[�����ϭl�v
 ����D�*�H��IOHk䄶RR�ϠM��Jk4i	�Ȑ�/�!1��#ΝA�l�g�XM�ݖ*���}6� �����/��n�����aš6DF �2 �/�JĊB���x�;�F��I 2��r��gl��w�hq�9Y�5;~�6�񻹘}������s2�7-,���=ϩ��u0V�#�Fw�c�N�,c{�ql�VF�tv��oDQ��qj��o��ͺ�j�uq���V�������}��ssN��E���ķĮ`=
%�ό��1���=
#�FFP�E�"�5�%����e�V6iܿ޼�mo���tB8xV@چ�Ù�j��􆚜D�(������K��`K� br���D��u2����;�7�r��sq�kC���1�.|Zr��c�tp��ǖW>Y쟌2��>5�&��C#mr�U���fƙ�Mnt���Y�ܸ-ʼg�Iw�B-�*�?�����'�z-[���8 L�b�S#���kv�\������:�g�t�u����l����?��#�[���t�E�<^���v�蒇DtX��J��a�!�u�B�X~�Ŀ�:Y��8x�>G�mp���p�R&T`�3:�B��Ӟ����;�io��a���0���$˰
~��c�mM���m�̳�U�;�ᣵ��sX2���(�˦��+RR� 1�Nm��;� ����	��o\Ì��C8���N[@JCw�`6�u6-q�t��6�z]V���	��4_�� R�_~ZH�0���LM
����?��>�Bl(���S ����Ǧ��h���)a���$˪P�	�����:���83N���[��2�O���'_oi��ՒTD����C@�Vn�ASŇ��"���.�ck�Uy��L���n�P�V�����P*�����r���v�1�Yˡ���>�3�Մg�Cs�lO9��sf�������QhN��fϹ���P�P�"�/���Pǝ+:���,j��+�A2�G�2���Ƴ��L��(GԂ�ГRpR&H��jBjdy"OK��vK u�d��mm�Q����8�9�F�d��}�{�of���;��P����Q��,J��q���2����
��#k�Ǔnb�݇�Eg֌8�8�bjV�F�\�n���P	��Eٱ�������F�3w;�l�����d��YR�uPІ,2~����`�@����ȅ���\͊���̫�3��]��'����r�d;ٞ��Z�i�G��s"��a
 �Fm�
�^W�Ns.y�[�;��U���cbP��!���$~^Y�&�|s0T�o���&�/sV�ɲ�R3e9)�Ԩ����N�8�&#�	W�1�.��!��%s�����9x�^�PVQjA�'��馆�3�6k���\�j��EZɶ�|���C���%WK�'��ɬr���K��y�_���r���s|5�#�A)�2!���5	�i�;U����4��R�]�R����Vd�^����m��~��_��(��v�9��`������t*�J(Hy��k�����t�X�����8����U�:	�j�`�8��LS|&)��RMi����F@\)J�E_�E��=���_�Ņ�$�	���>j����ٟ-��'8�������O~�G�p�ܓh�/��/)�d�
R��>[�q<B��ù8���?�G��	M�Yu7�--s������\o��*�-����F�i�;����9��V>Xƨ�C.��'�*0�O.�����$~w^Y��o��4�\��t.�1��̂�h8��p�2����㽒FpM*'c/�(\\��<v���J�p\^���w�� +٠�����Xw�=I��ⳟ\��c�[�1�a����'~∖Hb�ԡ�������<�9��#��ׯ��M�茉��a;��՟g[{~M�&�+fy��A�\��+�ͳr�浪�k9)S���M����k��e˺{��K>0=��<���Ϡp&h�
��L���J�w�Iih=x�4�r˗�����i��} w��2�vff8���q��X0�S��Z�E��aI��ß�q±V1D��c䀴�kh���1�9|�3�9�IH�c�A�A8�>�$�#���	�F�
��!}*z:Jk�RNP�.O�D��l����7�Vk����.����t���'�"��QF� �9R[�~�����{r.&*�I~�~C��ⰽ1w�(ը�q���f1~<K�;mHf�UZA�*�Nz,��m����IL6��	{-�<B]�P}����w�w����k���; �FIIYƃ�gL*ڷ�]2��O��1α�c��ˤ���w����H^���s��+�z-k��p
I-�ּ�9��Ԁ{���y:EM(� �4��Pe�0ǺK,@�Y�ɑ< }ҳ:�QKKm<�ޘ������[�*9λ%��2%Cǵڙf~�������~D� ���G �L�1��G]&�p.�e��yܗ�\Is�9:c�ύ�ВJ�t�j�Y���3lS۳NF��͘�\(<&�U~�S>��o�����Z�����*� K�S����.��v$�Y��EI�Ey������('�geC��s�F�A��	S��4M����-	&���~�`�4�k��s�A���:�z�5�Z�C2��.p�v+o�5��0����ukǩ�K:˱!�����*�z?�,A�E��������V���Nj��LJ���'>m�u/:E�b�7��k�YtrH��>Y6z�2v@���1�N��N��V�:�x���H���Ni =�H��1	�|D+v��jY���I���#��W�hz� �O�x���x����xԴ��2�;O�Im��ԨS�κ"��L�3z^��˒��6+7_W�������]��T�VaIM���*'^Ƹ��k _��%.x���Ό�'�Ho��7������\�O�o���E&c�0�:���8��PA��M�8���G\�8�D��ƩV0��� �1�P���t�5��L���>w,q�z-��'��I��*�OC`�����9�)x^���B�b�j�� �v�SJ �tw�����HW�{�3��g���4�l:�\rK3۹�z��<�ݥ\�l����E����OG�ٸnM��>H�8���`�[x��ɚ�hi��t�|���ef��	�p���s��UrA��v�Zc�T����F�{���fD%q�$@L;F��3� �"'5�V�-����w���^ku��U+���T�L�������2P�E��L�zQ�컼�3�OGlƆƘN�|���ZWY^���w�s���B. 0sE�2��2��4~��Oȅ�~�����N��'�����4���v��ݹ���{��r�nI[p	"�2/d�<WhӌyA��QIM�I�LS����� Nэ/��//�������'b�d]��$�Ok�KG+���ns��}?�>ۛ6��t��-��9�)��Pg��� ��D�	��������` R�/�K�3XX�X�l3\K]��JC$հ�$�w%��ꐷ\ 385�4��G ^e�
����ч����>�<A���@j DRK��p����XJG~Xm��E:-)�ia��-L���_�y$�`������K<<�s�g|�{�S
�[�tM�B��^Q"�S?�So��N_��'`��F��]�\�cn�mG�Ō����W��> 7[6�������/~IE���ښ� ��S����~����J�4 ���w$L)����%��/���{��	�����e�y�M7��r~�Yo�B�/9Ư=�ؒ�-Z�@8If�ġ-�R�Z����'�������>�nU:��j-hS����[/�d�ߵT�.Gj��P"�Y���5��x�L�I*$��y���~~������!iiy���Tº9ʱ�!衇J��ׯ}�k��ء�q
�K�x����QI�^�E|��F�7(@`���������e
A���x9 ���Z�A��r�8�[z�\}����>�SK�#;k��`�g����|тY�ȼa%�;���=/%��r?�Nxӛ�TJ(�n�V'�|_�_P��k
�9��l�U��xܛ�A}Q:ig��r�פ�>��?=R�����se�E�J$��=�yw_ϡk��ng�^fA8��4VDS�v�n���gc@q-��o��� X�TIJ����N�MP^j�`���v|$�'�@�@=��Z�H�@
C�Pm��pN�ǉ�%&A��oy�[�_��_+������%��X+0�(o� ,�E$�0Wğ���^���<P��^h�(��/��pٸ���&P)�1�+l;��M�Ox�S� n�$�x����Լ4{=�>�`���K�����<���/��/��|ei|�C�(���ȁ�N,�!��9�~k;^�nǤCE�L���8�a�����2#�`zd��r� �9��^k�h����\׺��,@[�<��Lzhk7H90��Eӂ3�,=�5�Z��:�2�;�65b?CR�^E{(*�akc�:��������ƨפ}��Ѐ�!N�3�s��{���s?�s��@��uH�� �@�{�mso����ŌfЄ/>:b>oG�Q;�ﴺa�y��>��E����������ұc\�������.Z-ׁw��0s`���W�������������u�5��ۿ��vr=���`�I��1�-�Ef1_,�Y����>��`���W�H��m�sZ¸]ہ����:h�<��a]�WϺ}ķW���x�+
 1���hY*lO��0��p��HWq�5@��K���\����1T/��T��	|x��_]ޑ9��7�qI�!���! �Ջe���i_��_ۼ��/l~��~�Ȃ��8ݠ `����Y U�2$�y(����;�8R�����^�L�I��:��p��Bf�<�'�q����bGs�Q-�FD�G��]�h(�;����
Au�4�4)���q�#��'I�tZ^���[�����ɖ�v��mM��l�hLLV)��t\�Wڅ�-��q�il�[/9�����4]M7	��0�|q�*][��W���	���F�6���^#�?3��Hϫ�jA�q���ь��]7G9������?+`
}/�jz�g�*v�Y�g��B�s��SN���P�xVh���������£#J�·jF�U���"X��qGd ӎ����P�<y9h	���
�'Z N3~%�/��\n��},��8�J���&��`�rq��g�.u0�q�d�����m�3=�I2�����dMm���{�+�fT���ٛ8'�r1��9�%��@���1� J�/�̾7�\^�qa8b��9�~g�U.� �1�>�4���u�k���ƍ�"�	��������jhj��,U�r��bA �Rp��4��d�{�myN~�b�9y/���vHŅ�΀W��^�aT��Թ���xM����vԍ�7�O���%R�/��/����� �أ!;8r[mX�I�ՄՍ�	��c�p��ꒋ1"������t�����!W��˭M��צ]���`�M��}��L+A 6D-���5���9�����x߭�:���e"��$����XT�
C>��`� � ���k��q�5���Z�
�s�I4�S��sƏ�w��~'���m�F�M�彩m̽P��`�u���=$yӥ}�
��O@5�����5�p�C:�td���� ��f�Z9D�ݳ\�&܎ǋŌ������%yHwS��r���ꏨ�f�$�J&�/�@W��x���vN;�ḁϲI���X��$�L��<Y���Y,��4j\�;��_?��hP���$t~~��T�`5�w�����$Ƿ��/����C��U\k��wU0��r��ߌy�_p�������,�c|y�t�^ř �o�����Q�Q$�)���D'�ǻ�.���,�/?mCA�6b�ءu�����}M���IR�`,%��Y+�Q��X0b��3�ɚ𸃠Yߐ��t��/6��4�SK�������CK`��R�v��0� ?9^���gpX�����zQ�Y�<��\�.,.����`)�.L(�52`~+�#u��N4�c�Ɋ���N��ܼ��� �J�;d�QFZ�^��#�d��?F�V�L�b�G 7�%�@��e�C�N�x�Q8(@��M�1�y3yV ؈��`��}w?��:-���W9@ՄYDT�2cϮ��Ԁs2Oǅm.qjM�ǒ�WV��<���e��ڹw��X� �+�����?���\��\���fŦ�����^aޖ`������,׋��]����}D:M�m�6t��5li'ʖ���6ʶC(/(
�UyWw#G��DH����43J&3��Y.|�Id4����^�4�|R�D�Pj��9��h���-�R���f�$�2��:�8(�����k��۾� ��~�����A��$�+��
O:@]��R��`�-�
�]��7:||<�`O��0�:h`�Q��R�e���f���������+��e_�A���(��� `��P3�s>˼yM�;Y䆙���&j�f��r�:<՘�����r+�+iN�4?1�	äo��˘Գ�Z�*mڟ'��B�T��7p?(�l	��?s���� -�3︟<�ڦ�8�7b��!��I�x��Fn�u��E%CF�K^����n��2��cwIg�JMǩH&Xg�"�[Z(����h���2�#�N؆��E01>����_:\4R��d;��A`�[�<�,�#�*�*�i�I=����Ⱥ�C4��PB�<����|6_:�)�����M�IN���{k	l���Em���(c葤ҩ�<I�J�	�1;�8s���"B>ǌ�F�.U�5��\���u��h�@F:��D����9o{��ʻ���>����P2���]��<3eP�W�+��j�$�����g�3��L:�J�?��c�D>���IZp�fzVYi�?�>�-�
���IEh��j�?�L~�!<0Vd��42���nI@�M�G�Nq�����=�@�=C��`�� �3������6�e�7z+�#�8a<耡cے�I���* ��;rHUf(�	[����w3+O��s&���q�Xs���*�������KA�����N\'�$܋g{��87���L�������,�����b�3D��YT�Ѩw��j�b6g�l'��h<-�0�>*3��?��J�����Y� )�j����rMz=��㚬pi�	@\�e/{Y�Q�F��Ȭ�Հ3f�,�W���������P��uO8���(��*���'��i�M[�3DK&)�4<J8�ag�(>g��%�̶�?����1����jق0���6��|��*@�ʔJV��Y;ƨ�\�|דD����zы^TƸad +��Q7Դ��-Fy�y~�s2輇�6-m��E�� '!�p�>r����k�	�%��N��� �>�����q�16.�A�`ry)_F�$7����А�wr�v*�!�y�k��C�;���0��?�S?�ܜ03��(M��e�y��̠2�Î7
BK��� 1aP�`�Y�t[�\Y�	�L^�P1��΅$-!�M�C[�\��Q�I��r[$5W~瘴l��� 67x徆�ɍf0�OJ�N�� ~9eD�.��8� �o��on|��bU�) 	�5�_���F� ^p<ֳ�������Z���%X��y�p�����͞A6J[��R:����L2L�O��Oj^��7ׯ�h>��?[�4���1�P**�����dU�=�Ƥb�����\)%G�Y��%7�xa;T�G�k3���@����9"�nQ��J��7*e�W�ˊ��N�\�5!�Y�G�8,`�NS��K���[���%#�$�o�"B,�W �����sė.�A�2 :��GY�s��	#�1p�`1GTPL쑣U[�Ӥ�zj��=�q���|S���Y  MFYB����u���
j�0������%>ڭ��ƿ뻾���;���e��1�F��rQ����,���r����Fb����5
^i�̦VM\����LZ�����a���d�����B�JY��O�����q`����6��%f���T&~�`��>v�&�⬐�X.iBls�r�i@;�lp}�\[���5��jIj5���8�@|���[��!���B��5r����A�t^�Y.�~�w�c�t�E"ǔ\*���sF$�J{dd��ajZ�|f�7c׹�U�)I�<+`��=�,
�S�V����=`���������u�ٗ���<�=�G#ϑ{?*�M�j��0�'�xtu�����_X^�	~%�Z ���Fc�Γ��@ ��uY�seup
�TMm��1���s@� �^�Z��Y������iz���j�i�aj���).Vj�75b@�j_��4uP'sMMX�~�1�Y_�- ���7���R���&�dn� ��s,�;[j�9�� H�$����AQ@Q�XY2V�_��Hh	C89��uZMe�IV#�|� �r�(��םj�<�s-B]��rĵr6�0���q����9��a�R���RM/�h~���<�h������bL��#Y�So,�Aʳf���������4�\Y�h��O��2����߮�6��(i�;Y��u�����Tn�%��EMg����E��4߭6|�Z`~F)V�m�X�:��R3<����  cq��q�?"˛r� z.�)�����e>����DI�5����\��ID%'��8�����7,'�����gý��wJ��1*-Fx���蘗�U�ח��y�CX��[k%�yoF3t�	�3q%�B��.��8�Y����W�Q_��o}�[�g�z�;%�Y�p��Sǂ�W��;��;CE\��m�d�K�!�J}7�h����!���?�>�1Ъ���-�!x� ߂��K�iMI�S��T�b_e���r,> �հDnnmeqr^�%�|�'�����ź��^�X3�6钌D�8Dʄ��[�%�㴐O9k�q,�<���:�sg񌭷x�A�0Ϩ�F`@�oJO��j����L�B*�=������7��1x;Tt��̧C
s�!ӱ�(A�����6��3�:�ģQ�D�z1��a���d�Ϡ�SNX��n ��q�vЛ�o8��9�,p#�ʨ���q�p�[	w���Ο�{ Tm13��.J-1N�qo|-�`h-�1�8�9f� (f���%c-w~q����_����n��c�z�'	mF���_���/��k[a��q���A8,�:X�?�EF����+�˱�k�$�������x|I!j8�\yv&}��^�sZ��+�������%����-���m9a���@q�M' �j�)ʧ���}�<8�L���Pc�����Lj5�h�	C?p�Zj�m+�c	��Nt���'����ݿ+��$p��4�jpy�:
�I�ǹ"`"����%�u9�,6��kX�Q�Z�>���~��o��r]�b���vQYWV�(Ƴ���F2�X ����S9�����` �)��iY�FP\��Yݝ�c���ɝfہ�������`r,A@U^�%M$�a!�& vb��� ���}�W�t��ۮ��b'Y@�Z�f5�����t&X��N�೚�C��{9RO��Y0�w�&
?L*�+�i�,��:�>S�SMm/�8X:�̮�Tz ��,c�}7��3��g��vN�$�/Ǡ�RF�9XN闬֦��u,�mq�,��s/J�I�A*ù�iھc.��8�xN��N��y� �Ĺ.��nz��>IRz9��,a�������&�ф�����軓%#4L�*9?8q&�+sZ��[�X3��)�#ﵕ��U���p�Ϛ��@k�&�"�R���C�{�/%?�|5O�RƔuX�_��{�Np�P�E�c�C�;D�X�`O��Ys�1��o�[`F?����*`f�|i��'��nV����\VY'��(�ssQƣҿ�ч�H���uWb�b�fQ��j��R#1[��;�ZD������V.Oj�A����c�!�t@��zr��
��HM1��R4�����ȥ��G����s�i��ؤ�q�=�������1ƽ���:M8ۢ�<\���(�~�����*�Z��(e��C��ƹ�dg��]܆9�(N&$'nz�kn�E*M�Ui+�:�A�OXT-5��H�B�֨\p9�T����:,��@̤���\�	��Ka��
�z�9�D6�Y�T�ۈ	�I� ZgY;Bz�{?���=�(-��Ƽ��P����2��q�^����c�&�n��� ��C~M�;�6�E�9�
�#F�j@��A=8�<�֞��VҏwI���-��c�41iUHZ�u�0 9F�u,���Z�TcG�㽾��ݑ[N@�FEj�n��C�{fVYf�%���]8�gH��\f�'�h�7���n.�g�� ������p �5���w; #�N�Bm�d�4�2?�ZH=�:u+�'�8F�'1�>�`� ������4r�[6��u#�w��Aҁ��?������+_j"�[()?ñ�ְP�Mm^P`��z�e(NIH���+�
�Wq��%�h�+5�Kq̝Vj �H�U���� ��Ť�T3�����ñ`VyJsP�N���H�' KG���/^�n����yV�c� sg�?�O���cܬ�5��rH��2�<���&/�q(S��2ؑ?MFk��*,�`|�r"/f�3��EM��#��}�� �`��"߭�b�tC��sn����\�V.WrqK>���2��H�7����ke�ǆ�R֞6�غ���9��v�����@VU�y�ȵ������PM'��s�C�;<6kN��:���JXu�Eʺ{]�p2O��-屲�1w)�d]U3�6	q��r<mb&��5�g�{��I�d�a2�I�)�U�����L��&��ˑ$
?#q���n�Ԥj�Q�5ـ1a�+=���6���ƕ#��qh��,Uh�E�.˙����sezr��Ҏ�t̩A�I���6$�$	������Eh_\4W|�ս
����6�4�ɸ%A�d������ Ð%wp���.��z@Mذd��9 WZ��U$�]}X/}�KK}
��	��Q�p��ʽ�61UD�\���ǥ*0m>��NI��o���/��|�V�c�=L�ɰC��^S.?7�o&��l�1`�	7�x����W�$������L4��*O|����
�l�U�;�l�[��)�Ǜ�f+گގ�	1?2Hm��'Z����~�k���e�;�ȝ5���*�H֡ �~��8���F�P��1@d�7��:/���;e >��3�[R���D��hՀ�:��G>�4qd�L�����_��R���g����4,/kf : 3�ٍM]��/]h<��f�fX 2��u�S+'���h����P���O*{��5ݐ�+]��s�� �i$�kG�O.� 3���Ea���u�+;�ґ=d�x�[����/�r���^��ׅ�$Ȩ]��ec��z�q�wX��k��֯�t���B�!�@�?���`��SǍ��u�Xx��q9���t�w$����K�dD��R�H�wr�逳�+0�u��3N��05A�k�E���o*9�Z�!o\�qc��J�*m�~G��̴h��X���:�d|��D]bv�aAr/F�CF����h�:2"(�Z����Va��#(4�3�E���g6�IJ�~PЄ��O�ce-'|p���C��bC��i�Xn<�	���E�ç��{�!��f��"/(�MU#4ƕdg�׽���m���7ӎ�B����z�j�j_f��~x�x�+W�݌;���f��3lĸj+��+y�ޔmۣ!Grq��j<��I�k���A.F\ۺ���1���ܚP.Y�$(�=���M�w�x,��ϡ{T�=��I;��G�8�������~��e����sj��t3O~������Sk6�LcK�q�x�(�`��;�V�����U�Z.����)�j)��\��I~����!������&Ub�r_+�Y����(�jÙ�9��9��h�`T�Q'ֳ��;��-�OGts����ޛ ݚ������t��!	�$l@.*�6(� �BDEL0�������[7Cݾ7�R�U^��X
j;&�hd0� *�DTEiA���3|�������o�o�=������~N���;�w�g=���4G���p���zsn8F�W��k��?�K(A��X�Y7t�L�=��O.������d�������Jg�@�T0�w�wO�Uy���������'��Ex�x0��d���K�����;��5��N�����e�s���>��W�bȓ����U��f��z����1��l

Q��I��@�Ș�$NA��~-�35�ǲ�����4�=X��]=#��X5'4��Ve�-��1WT�E�u�Y��H55�� (��/(�A��>P4V�Vf��#���ۻ�����\���F��3�)�ڎ)��Iyű�#_��fO^�A�7���V��؊��1l�]+|{���]5ƶ�b7�J����]߮&�����
�-E��*B�΢H;��f��#`r�z���������A�n��Ğ���G
l����,���:LT�Z�(�ۋ
���},�a��� '�,���9�sk��	 *��6M���gx	d?���}'Ha4�Co|��LD��r��,T�"� "�GU�fi[�E� f������e�Ls���-���w����.|��r,fgϻl��EH^\ೡ8�Af .+; ��gb�a�j��;M��	��K_�Ҳ8P������9���;4@�Ƚ ����<es�v-^z�$̆vk��\3������U�yl��O�y11�r���b��J�<�iO+*�z���7�,��t������j����z�"J�ű����ѽ�6�s,�@#[S{�^i:��À�.��%���/��0�j+2L���l���,lT;N�=��)@E�u��h�`L'�0��Ƈ�Fd���J�4�\L���	M��/���b�ӱ�=,��o�!� *���Y#�%5q%��Gi�RXr����q�(#ҙ����؏��t�2�r�P��"�ǋE�?�ma�f�/��S����l�rL�*�jM�j��J-s�$�4c�b���Y���ۄWV����䳞�����|�����:|�Cz@>,� A���Z�0P_�Aa"S�=+X�V
M�"��U*�c��(Tā��3)���p���8�m�'kH�����Z1�d��DӪt��չ`m��D�h�n#L���X�H��qW%�}����2OL�}���Mۅ�f|ޮ1n�c�b0�>_ބ BK��.+�ȍ?%~��$���c��Sё����4K�\�	�Z���s�8�M^�M��z1�o��V�	��	p�����s\{�E�
�D���at�&M}B���Q��R�L�{j.�A8͟���*��h�����q��Ak뭀�:?U�VWNs+jB�����<���p���8�`x7yP���v�+�+���EG�h�߻�S��.�t`���p�����k��%ӯ��������ӎ�;s�3�4md�����N ��ԩQ,zv�B4Mc���d�h��plB�9ǋ��mn���ow[��s\��"�[�h���X���7���T��N��b�SV�ct�)ɂ��ղ��(@�����\,f9���{k�P�z~֙�3tK\�g���6^�;}'�d�ۜA�~�`l����9��W���1��M{��z���]d��L2���� �)~�l�y�D;	���Eă�UV$�icU�h��u؉X�AԬv"?����HWAC�M������P��`�9��Ύ[*Mz�8��w�h6�S����6���ȏt��#���R�K�㱪��&B��$�c�H��`Z�k|��O?�я)����G�3���w��	�V���y�4���`�$�D_��ѧL
����3�!U\7.�f�H���q�F��lc"�4�-
�����n
8�4NI�.���~��F,��\�}&����U`:O���D:�;�09�w���Y<�ߐ+h�FY]��-����b�����ћ#�M����Fsթ�J�/�ˆ�A8�0d�Y�B�blN<��AxX&:Bt�Ȥ�qH�
����Y��o,�@��6�;��`:�cJa�6VQ��ɐ����n�v���X�j�B�	��� ��Ƞ�2ݽ��6�K^P�.�BȀ���n�i�;K��RMN�h��Z�g�i�7:22I�K��+_���=�cxG�Y_8��y��w�}�k���'�3�k!;@�P�\h>�}Ӂσ�%��q�]�V��'���:��3g�96���7G��PV����0l�P�����I�]疓8�aVI2X�ϱf:����0
B��;�u��7xn�3z\���H!4�j[e���.s��Y�=��7��Z}��L��|��2���e�l�{��a,�w�Z�?*���U�y-2��^���ٽ��,��DE���U���dY�}���s�}mҪ���~�g�h�|���F�#7�]6?�!@��_�C�r��aH��A �!�-��R�4|-ې�ؤ�L�0��(/�ى�2�'�^���5��/W#+si۲��0P������k�f�'I���Y:��/��0�����ogz�3����"���6�Ӆ	�&�&�D���03Q�N(��wm˽u>�6@������~� Nހ@�?�3?S�Ђ��L�:��� d@��K��<^I�\����F�K?DF������4e���]3ID��?����<��uו�c�E>`�@&������a��)� M���KS��nD���1��ʨ�9*�\Ͷ7�J�'�c*U ;6���������]>���-���(��,�j��ʢ#�Wņs�_���j$�E�μk؍�&�"X����*���1��ܓ�g˶�*}�_�2��q;w�t2�L7�dL��ݰ*�h[�\���X5��`a4"���P��K]LˮwP��E���F�(�(�^��-� ���_��.�i��o~sɠ���^f�M��Yo�vQ��v��?�M~��ʶQ�	�-�0�o��n���ډ�����X��)ҭ�R�@Ⱥ��!%; ��9�/� ����-E���5(;���=(�=���U�h��L0��Ô|�Ȕ夽h�_� ��hpb����#4��H��Ʋ�4Ҍ�=��@''<���U ��(���p=
azR�e�C��W���{��	c�	�z���9 ���E-�23
�N����N��R}+�Vy?*e���y,�	��[y�o4��&̱A<��
z�賙v~�'ծ���F{M�W.O{&�p����;G��_򒗔�#I���
��J�o4��{��.�S3��(�8N���R��a9��ن����k%�l<����`�C��횒2���?H�4�X-0���B�������B蘧V�� ��\�UuI8�įx�+J�Z��܃,6��sMl�fM��g�d��R�T���e��<�����i��-�뭴S��s��h0NW�;n�� .T_���<NQZ�M%�	������d����
c�;�!���U��&ev��?���k�gr�D<���7���\���f����na�<�ϻ�գ�������6����A<&� �Ǥ�Y�E�E6�Y8�M�����"G5fA���Y&�M�RF�)�c��(:�ع��}�|o�">�o� ������S�f�c�MԨ�>��h��r��-S0�{���)LxV�k����*�u�ݍ�zt �T��P�l�"4B�����<k��,B8kxʼzD�CN�ݝ׻ݽL�2���T���.�%]qFB�餃���R�jgdڻ�}����{������S%�����{
�#�����׷��嶟7'����v���+��~�n���"�����#$U�4���Ѱ���D���0���|�)�L�wz�H��KAݠ �j��5@q��F3�<�U��V������=�3�B��I&�B4lL���BK��6i �}S��i�0s�e>����~�b�G�^Ď�G,�� 1�Fަ��o�����^]�e��n��]�J�C�)@e����O��v�Q��ʫGgPro+�$�ێ��(�S�;.��i��e-{��8�����O�Y��/�՞k��2�D3��&v����,��A���pVPf�}��ש�h��qg��eV�jw�I!��f�x�W:��\h��wF,��E�y�����6��5�<��ܡ���%h�nLR��c�U#\���>��	��w�q�c�&�c*g��>Xm����J�i�I;��"4���ͫKt�g>�?�9�
ܜ��e`�D0�v>����ʕ��_��W��=n��꫋�x\Rs�tG�F��%]W�㤌M���z@��5�J�c�C�6��s�E�{Ht��̅ӱ��@�z�T��m�ud��, q^���] 8�{��ģ�a������ݑ]8D��v��6-+#ۅ����e/+�e����E%���!J���[M���S��a�G�Z���1�����\��SI�Y��-����	S�b�5��}a�6Cm�G=��%n���G�:�!�>(�/B�L94ˊ�	"���H���/.i�=&>uEA�T�'F�X�D����b��B���b��R���ksE�zҧ��ʦ��k�v^�7mf��QL��;�%师L�]O&�1� [�Y���A|�pD�����^�c�
�y�!� ��Q(���zU�D�Tl$s��0)�.L��Fq��F1�,N$?�W���V�>چ�=���1�R$��}��G�?�%������kvw� te�\�3Ep"����q�dh��"�R�[��L
%�9�)��r�������X�7��=>򑏔�,jU���U�z���/�ʖH�Kq���:k.B�ƐH �U��y��[� ��S�{��Jb-�=f��� $*��|Ϝ�t���"!� cY+�ۨ@��A|F���r<s�v�2]��y�5��(ؤ����,��M�Bc��_����D*f�c���e)Y�� %� SBa�[@����枤]�<�?�pݤc��6Gee�N��-%yb�D��続�?���.� 0B�,��at����A ����P'&�c�Q\����F3MWۙ�<M![hCU]�]�N�z��C0k�f5�bW���/m}�������B)l�SC����S�0�R�[)��ַ���[��"8���7�s$Z���b^q-�^��W4��?���LJ-�Ë\��o�!��;���M<>�������Y�/��/ԙ6�����ۿ�|�h �gĉfv-u"xVk##{�~]�X����h���g���ݐNw�D�`�@�q|ڝ��I+���Bx@�Q���&�s�O�6��qkY]>��/��-x8:,��
F��3�nR�v�D��M���6��Yp�O�QR�J�!C_L�>���ժ��n.�.�D����t%W}��R�Hdz�k��R�?�)�cjB9���5���(��Nt��f�|��8�����qJY��y��h�F"���\�hv@����|���)�!�)"Rw�ܛ>@���2������E�z�օ����	��Dv�!�耢s#T�5`���?C�l�Q��R	E�ⲫRЮ(%�u��Xcu����&HT%��4�cݞ����!H�ņ�I��G��o��b��ZT]���<P�5�3U9=��t|����"��v^��MӁ�c��^���)8�n��v>� S-t�o���`3��cR�}
��Qȝ!8�H�x�32�4��_CHQ�-t�-���)�W�)�ۍJ��`����h�����o�뻾��0i�*h8ܨ��%s��ұ�9}�s#G �`)���	�J<2�_���Q.����uD.��)��;�wW��JO�����>����ǉ��|i0O�J���5�#��]��0��~闦�`Z0^���A]�� ~ғ�����e�����#�fy�Y�e����<���y�9�	y�Ь~��T��\����'��K�~J6��o,��Ŝ�0��O����
#��bYF�ٽ�mo+�F��s 4�!,�� &:	r;M�鼭�$�W����q�")ʠt"" _f�������E����W�(R(sM^,PԞ�gʫ4:N.��$q�M�m;�:4LIU��ϕ���;褁�(��Ƴ	��0M���5�3�-��=�N�qڮ.��㦋�?���q��(h��;�EW"*�~���A�|��v;,�55ZH�� "~V�[{49��
A�����s�"D�%�a�-��=�g��X� j�̡4�%R�G
մ'_u1��1���_�j�T?P�	j�g�.���!Wڬ��a���bǪf�}t_�e������A����Ԁ&6e&�d���:�B4�ݗ��<Um���&�r5)�Paw��8�.K�b�l%�ˍ&2�Ӆ#�\��ϟ}��jW�h\J�w�!j[$ktk����O��X�+�fP��v��-��l��KA C��^��-37,b�KI_L��]�W��2�%��Ō�v�d�vv��������B=A���v�"h� �xf[iFМ��]��,@�%§>gdM�}ҡ��X�tGw�#g��hj0�]5��l��kj�I�Ţ�1��y�����h�B�`8�ť,����K���N쬧��s"c`u��(��03���:�����/�1<NT�����~�4�t5W%�ۧ�}�E�9zs���7��|)�0i����Jngb�_���6���Rt�]�4ϔ��|'�~���(��b/���rG���6�4a�Ӟ�'�iF�(�t �����^�"��xv���6k�'�%Q���ފ��޽9��"�Xf)�NR��;�	���g�-�� ]�,5̀�&��6;S�+�)�y�ܺ��i���,9�ߏ�v���*�j&�E[�_��[�id�k
_��)��T�S0�7?�"\�s4�n����s��m�o�t%"�p"Z�1�t%��e�>Ʌ� ��h�Vi�Җ���b�j�U#�e���J���,�(9���P�}��"T���lQ�z��E��������4�=}�������v�&2�kߏ)[��L6��!��<��|�WVS�f�-Qs��t�mH�q�/�ڶ3^W3�Ϻh�̣4�@�5_��OZ,�WT)n��q�6�>&�?*�i< �_j�[���ߙ5��VЋ��൬qꠤ�@�D4mx/�;Zd��g��8��g��Y���^S�Y?�(��e�Mڹ4٤-�g�g��يI�?���z��皕U���lm����W����LP�p,�{�>����e։��&e[D0�(������E��ϑ߉^�l��\�����Tצ��Od%�QH;o�
��i�NԘť<5/�R0j�����z{�4Zx=3�fQ �u|'�)��I>���=����{Q~���_.^8#{T���vA�H�[��Wzڋ�9e��B�n�p��z�R
�X(���T-j�!c�ex�� ��n�ݐ�\]�1�M2�� ��|�'���>��ƿm�!��iCS�7�s��u?���S8���A�/��E�6u2ʇ�s�ZX���m�hš���W�Q�G5n���J��r��v{啋���>S�]���9n�	B���N2R��%:�{��˩ۚ�L�C�Q^�k������	`��5���;���9g�f���U)s��Hj��>9��h08}�Hx8,����7L����[ؘ�v�^Yo��<;����J�ꖅ�U?\��xu:"�.Ls�/��m��-J�W`��9	jЫ<��|�(�A��\��������&k�f��j��j�,sRM�A��XMl+��^iphǃ�����N����ś����]^@�����~l,P��]�{������X�
9�,�(���@�xU���Җ��+?�b��Zjx)�Ҷ�ɝB@��e&��Ț���r#%��!�Ŧ(�y��ㇿ/���K�M��a)ۂ�^q�Q�#VVze��7��;U���W}�_o�k;��&ج�.i���$ۇL��C.0,F��6��w�@�E��*`S��d*�tl'����v�ʩ��DE
�p�B@�L�oE6�(�>�������!(0 �ͧ��\�Y⹇��t۰�V~����?�R�����0��֊ݝ�V����F�=��U� �[�M�sͥL���!��妗YQ�1��4�ɳ�δv�e�	XD5*�-j�^���IJ��m�Z�M>��q0o���0m�|��q�k�igتQ�>���"?i����]r	\S�%t����n��6���\!|������ŧ�����`�ln��'ڎm;���}�U͉S��yV��<�9�f�<t.e�O�5m�LΧCefW>�w����&�H�"�v���
X3�,b�03���J�n�"�SX/r�uۇ��b���R�+>��`d�Y2Q����.D�`/��������+��x��;K��,��u��w��޻]�A���ܫ���-2�a�p��=�����j+�vn�N4���#�B�����Љ>3�_��9���=c��
�=��%: �(�+�T@��m���C~OM��E�lw�-��kB���q�N�癙�TP�w�#Jfo��������������<��>�*(mY�X0�w��m�7ƍl��6�Q�_��<�1k�[t<<� _8Q�	a����.#(`�,jz�K�j߻�xgb�U��	��YE�Gu&��QϘB*2}
&'N2,��
��#���
T�B�.
]�*��Q��1��S��~�{��ez��B.l/%R�kʊ�ET���b۝h1�Z}p~��Э�쵼�}��f�s�����M�$x~����Ѣ�m&H�]p7N5�'O7ۣ����[��k>��ϵ���| \��=6��x��V���Xi�<��$66P�q�P"N����3�{�
�ź��l��`'�� IW�RX�9���k��e��A�Tf��o���ϥ�'���Ԗ��0s��6��ŏc�1���񿌜?��~��T�a�i�>��n��{p�w~k\�z��fY�9|�ӓݖ�'.�6P��qX���2��}m)pMiL�����z���m�D�aJ��d*���믟�.�`��&U�e�d:J���aS4��ך�]a;&&��|��3,C�&�'��?���/E�a������l�����Ye>� �F�w�£��o�Fi�y�9gx��XG��h�;c4ǳ=�Y�5�}̣���<Ӝ���f������|��vY�G���k����<�-��ۅ���͕ts~�b���{��8�΢a�x��#�wߗ��Z��@�0ο����h��O�Q����UĘ����}�X5����$+d���2������ȗ*f�����t�97�'�!��[��N�;0��^(��s�1��1�L~��~m��5�����/x��_��_�.|o��Tx��	��w(�A.���XC���:����$�7 �Iz�t�R�m���fj��n��mM����*���vyQ���(�/�R��~��`wh�ߩJa:����#�!9��� 08���9�( �+Ì8a�hv೓���A@�L��炥���h#��>����	R�fҊ��x�ϳe�	߻ןU��M��`� Y_�Ew�B�h�h�qeԎI�]�Ϸm�Ex�9��;����~�X�&�/-/��yT�4W�n5""�'�����>����~\�ܱ}�U�K�PD?#���'~�B9�w���uP��)���.�C�]6~jc���F�}���@Q�����f��1i�E�r'�e��|�3�Yd�;����ۿ���w�/�����R_�
6�Q��� y�<�AQ�S��]�R�����q-�sG�]I��+��3�	l������U$��oM
2��ЎRhhc���F�S:�� ��R�w����=�!�(�e�e��e�P�Iv%��%�禭++Q�7���P6h�E��̕i�Y�U��Z��2��6hW��z�3�'×�3ĉ��]sU���'�5�|Xkm[��^iE�U����볛줟v������jy�-kZ����Ҿ�a1b<W[�^8-�w`E�h��t>��4U�4�i6s.��N��hU��ڝN;�N!�b������W'sn�OĶ��&�;��ֺ���3"@���}��1���d$��Hǝ���h~q~z_��fJ�6#Tv��H�3��#O[n[�>̰���ꇚ��E��Uk̼�J� )&2���k�����!|Q�0=`�0�	"�2���_�I��P�.yL�<2�q�m��O鑌b�8�hXz�N����.���ҟ8i'כ>߰��J�ƈ05�o���$��L�a	^[��V���7�9�(o��֬�֊ѡ]^�Ai'�N�R�BL���s����"�ü�ͻw��-z�}7���X?�A��&�Ź�%��g47�tS�� &���1̽Պ]8�؇i��|�L��ҾX����eqWO6����9���
��z�)�^�$�r���s��PG� _lS\��VɬF%Cw1�/��y�<k����x�.�K{�I��Ьg�eJ�O
�����c43�tǉ�@Л��p,C�G�yI�W���N�a˞8��Rk�j��o����kMo@��N9��|�R
�Y<Q/�)h��Z�5�ݳ�"_��˜�ۜ'���e���_��c��� bh��ԴhLp�y�F���%K�*�5A�#�Y=��w@���	�ֶi騿���J8��r����)��N�C�U���i��A�a�����a�bl�f�m������l���`L�搮����Yh �LM�PD����:��eֽ�����i���f֯{df9h��[e��qZ��>�Zi�ޤ��j:����M����iX5ū5u�y쬿��,�t��� ��E/zQ�z	���# eK���ۈ�S����V�7��SKT �N��W����	���m��6ڝ�{mD�x�4U/8�g���C��ԙ75z� ^�4�{U�/�t�0�N�����jd�Up�Z�}���,4=��௙d����H��5tI�x��X}�.ҽ&�����V�)O�����D�p��¼ԗh�3�r~����y��^�ۼEt���K�*H�-5�8�)�&M	_�5_Ӽ��/-�  b^D��	�_����#������n��פ?'�(iZ��Fo�=�Ӗ{��c����	��1.�	Qgޘ.;�Q����ˈ�!�9Z����f����P�e4O��b�Y���N�E(��e�E��^`�۾���wfo�%�gԢ��T�����7,/2��ʫ!ss�����lM�d�]d��Z4��T�zQ��w�~�Z�C�JS�֏��-�B����w��(ur��~���9S��h�ܹP�����g��&�ű<L�+�}���s7����(-3�߆�X�^��f���?�8�D�؀�|��ߘ#>��UE�'g�X������y��"J�j}�A�<�;o�^��R#�"�g&�C��{�S�ؤ05[n����1KfX�p�����^��V����������fH�ۨ���K�,1�O�� ϲ)׿մ/Mf����z�����"��:l�K�/1�8�	�\��FL�<�D��g����6�/J�Ub��Od�>ZieоW��!j[#�sDz�w� �{P���}u���N�'RP�@)<�	OxBY�f�5�H�
Z,Ę��؂Q-�jA�`�+���v�SK����M��,;aݧyݬv������f\%m�B[��vnvz�6��IXk��m��ˠ�v|G؁����Aqᵂ�x��乊�btI��y�z�f�f�2�s�WW�ټs�^��j��"g�aH�W�V�ٝ�цMK�j��Y�7?ב^�-A_��P;X_/��hF��[��k�hgP�K]����n��������N�ґ����<xE?�яN�T���h��l v�uQY�}��t�����p��k���.2o� �>�'>��0YM���MR=i�Y��@0"ǳ �����$b��}�q��CaWs��ZG۹^��ELX&NТ崇�w���������4=ܭ3������I2�,�h֦��JU��n=��K������,B����nF�ԞX/μ��|s)Q-h�����^�ѵ�^;�D˰Ay��C�E����HL�ٝ!�y�i�R ��[��LQ�ݐ�=$V�v��;"H�'Z(�Ȑ��t�{lF8��7��M���}�ו�A��[��ɟ��TF�j�L�x5S�
]�ߝ�Y���`YQmy5ҬA��"��m_���<ٮ<��q��k�d3ȇ�F�j���|utD��f�H��2��!� S:�2�54�/"S�3�;�b�
�4�X��A�ٸ�����r-�d�Qf%���j2EڊP�Ǆ�/h/��xle,Rz�y7>۾6������2,}ɤ�=��Q]����λJ�Й��������R:mP��JɐM"ن�D1F�8���x` o�dʵ-/�E>W�n?���<ِ�����U^Ÿ�Y���"���k����M�y�{
����y��)r2[sY�h�\��0��3��̴�+�%1�+��υެIgh����xf��E�u�����2��H) $m�ޟ��N]ն_HЗ�X����3( �e�����j�S@%��]]�(+�)���+2��+M>H2]�\|�������䋿��(G�xP(�Zv���(p���I]�9 ��5r G+�Y�r7[&�s����X��s]�|��y�4���l{d�=���n}�G��eә�w˜.E��Z�{w��8q� tn�m��z���N��7�����Qn�4��(�jd�����V��O�������wi��t�V�V�B���|+�g55���u(HL1���� \��1V�Ԅh�*yV��!�3Y["͌������z�)/إb	��h��}�@�� ���y�\uQ}�D��!�.�q�K�Ej3i2��)��W�H�5���T@)� �m�D�(�G[M����N��_��_++*�"H� k�9�yN�Mj���R͟g���Y����Ⓕ�tY�&pPUwl{�^�k��.��R�rR��<�h��dz�5�p���_�+�n=�]���¤��2<�2�^,'Ka����8�����]dW6�;eLh\Vxe|͉íe�r�������M�Hr�X�9��7x������-:͚�FiG�R4�9e��B�ڿ��碑%S}>�Mm�9#R��ѥ�ڛ���"�5�P��ڃ %�־2?WP.H�P�P�Unh�Ȩ�Lh�����G���##��X��j�LS�A�DW�0�Z��&U�\� V>�T���&��*`�O��OM;S��E g�@D���m��Y��L&�h�{�*��".�q�r��$�x�h)LHg��c�J�QSH:I�N.�9�]h{��Y��[��!@���9�i���}�k]�jd|pE��q���cĿ3�)��z�_x�QmW;�+�Π�#��X�{���1�P�k֡�"��p�:s̶["��t5{h*��꼁rA�9D�]���	��^����������� P[��L���vhb��n��g�1���[�ȹ�};�~�GG,�'�������1v���f��Pm�H�,�a�h��a����ud�h��1g�2I��b���� ��i���\]s���Y�G���+�ղ�}:gr��{:F]XH(H�
�<�����a_om�0���ń��.D�����N�s4A�͸�Ψ��Y)���NwS.qÍN`�ž��#�7�C$/U��1�Ij�R�Q�m*D)e��X���s�\�e���^���ҧ /��9�����b߅�g�,�Bʸr�����e1b�	J��T#��o�ʚ	�j9������ZDN�;�>M��Gp��ϊs枳�����!'u2\��$(䤭O(��iO{ZA��z���+��+eP�v�����"��,]�=;�P��D�P)�Dz����<GT�0�ڳ��(;M	N��;�6gU,��ue�e��_
���{��p~���Z|�GeM�h�����[�IGc�:�.�}څ}�Ef��˽
���/e�ܔ��r�M;����B�6��p�N�.�s-CN�Ye{�.��{��N�E�<��gKg|���[%��p��/������r�Y���H$#"DЖ��<��!yuTJ��4�j���R�M�x�����4L롧�*Q�<���D߭˩
��4C;\]DPt\����o
9��5�)�'���Q,ЬP��j��^D�z��hK�p4�v-��
�I�v��L�k���Q;B��H���P��
�,l�ئF�t�jt�n�����-���&��m���λ2�<2�t��h��>z&5��?�-�A���d�	�V�����p�Slė2�����^�M>5N�hj��0�\�S8v	QH�r>A�O��(��U(�춋߻ڂ%����8��TL�:|F;��>�k��v>EE�ڴ���9� ��s��B�y��_�d����V%Ul/͸�֢sk��O5�U<U�o{�ۊ�Fx;6=�ڗ��t��b��	�����g���:���~I���T��ez�#QWmk��� �h�n�����=�jh��`l<�d�L�kT�.x�q�[���k������@a-�^�p8�y��F��C�u,뱆R t
�м�R�L�ؕ�=�G�]>��8�H�D��x�͋_���)OyJq�s?�I�"��L:�dSon���<LԿ������s�S[8u@�fd����P"Vn�=�F����Fꕖ�~��)�)[���
_h?��yt���4N�m���w&;p7:�,ҥ,όZ����[�����y Ӽ���E�%�XcзU��ַ�=X���B@S_BP!�U�.k�祶�5 ��4y֣������R�ⶻok>��6w������Ul>�'٬�Ϫ�:�h�����I5�T�ۢ�v9��J��$����E�y�7)��w���σ}�t5J�t�u����O� �2���1�"{��V�yx�m�]4��}i��j�Ӷ�誨IS'*�*1�S(���^�2J�b~.��Y��B\M��y�Zi��4£�e��Y����2�Nc��[�~6��vK�ܼ�&�M��_p�K�q9�aA�<��z]A�~�|
[Mځ1I�����S����e�i�ά`���#��hsí�R�l�����D8����T���p�ݦ�Xt��6v�N �ź���ric,���܅�b�OA�^�+��f�ʌ���[o4�s�pυ�.�t,�5^|-q�r��dw�@�Z���!�4h##������y������<� ϸ���7*��iW��v��}���-��<��YIw��������OpW�e�?,]�4)�>�É����5��񽴷�����l�w����d��y�(��D���0��Q[v���0��cȘk��m���a��/'�?Zj�Xf�Q���X?Lx0KlV��A���Mx4)��Oa8�3�F��E,8�i�o���qͯ��U�ƌU��+
�Ġ�@9bA۠��ݬ���e�_:�2���zj�I��7��w���dS�f����]F��r�ڬ�+�n�E+Ee�V]Z�;�����-ȳ��kHa�M9ߧ��Aa|�tX��7��㘳��ڂ35�cY��ΰ>� �L��GQ�0��u�	K�LQ�暃N��)�ks��ze:m쾬��ԟ\�ܹ#�,cc?!��(6b=ތ	������'��~�p����3��#��a�'�2S���2� ʪ���'�����[D�c�"[^#�-b5��a͸�	#�<��7M8˦��	SE�Wb�.�8 ����/~�#�����N�$�R�	 �;�9䠂q�����A:
JA��m��2�明<K�@"E�נ�eg�Y�59�FK�#.'��z��)#Q"�6�E��2�3ge���A��I�>�@��d�Q��F³4;�`���s�w\����1��e:�h� �}�0�=Z
s�tJ֛H�|�s҃t_P��*!@��=�n�iɐZ��Y��g8��i�.{!��D�ڈ�,6ߥԤY8�����R����Z$�����dĒ����^��xt�s�q9�"a8�zT�.C�VĂ��fM��`�ti�|�++�e�4=d�nskqw��A��Lz����.{$�l�3��(���YK�e�N]�X�=��=H� ��-k��)3T�4�oC�F mpt��� �G���W����]֮XF2��8m�҃t�R]WSD�,�G��eM�4A̪i�`��^��0dQlw� �(�y�Ö���j5~�#�K��N�3�򸖉%x��u7ǝw
O�@O��-�Q1�1�n��*b�Z�Z,��?큦�&:�Tt%vͦ&+�s���O�B�X���7E��	kvXa�ο�[.����g=�\볟�ly���}��ԧ�xn§���չ��Zͼ~��G���_��e�6�~��X�Q'+�j}A����ig��ǔ�F�pj���Ju2�	[1�0�e]����u���S@]A�߅��~���wwW�L�L��N��v��`K��
���3
����������˱0E���暹����~��C�^L�����^َ�Ҝ#c~��/��	QGR�H���]OO'�&]����~i/�X��)�ԏ|�#�lN8ⴟ���6Ox���}�c�w~s�F������2&��{�W���r_V6d�~�~�,z*�]�X�RO��E���GuD@�-vM4�Lهf�AY;���4#~��`,��a����yO���l/�.6|����y�K_zA�^H��w��쀮V�M��Me�,��q�-6�u�u��L1���C<:�I��")�f 	1��l�����&�Գ�W�Y<\�Gx���!L�!��gU~h�������w�5KU��qYr�@(���-8��)w�6�ߝ�3��c���*Z���,��g��1���?��JSR]�oY�.�ܭ7�??/"3��_7��><�a�5��nj����<7�����٘<�n-��b��\lsOC��eȚg���u��a�������i�^���ovmI�0*C��=���뻦��D�	  ��8��H$��=*r?����]�2!�dr��
=�e��d`�8N
�Da�f���@��x+jy}���+�Nn��/����_�����Yί$c�	'��.�ۏ��$"�V0��\Y�hrh�ews�r�pr��Yu�_}��g?{�N���N�c*J�T����+['���~�Y�A`$�U[��� wa�w�Ff�~��8��b�
(�͢e��V��q8�D��s?�Ð��>5:$N����~N��W�m�|ge=?���^J����C�9����sKV���r3�.�F"}�e�p����	z���wP�{�s]l�hkɷ���P�U�Ml���]��1���D�����`��,b���P�P��-����?��He����-������� ew
8(��JN�܄�3��}��Y^�.H���18�D��#%���z��D�j	)DT�sgm�:n�Fѹ�0��6z>�0�dͣY}4K��f�Ft	�d|<^j�ٮ�C~ss^(5�	G����l����D���D�:��oc��un^+�v��[d�耓���2�L�JS���c-]{g��9T�at��ǧ�`2!�q�bR}��xGE6��N[0�0�Cާ����� Ƴ�Șŏ������|���k�A�v�5�R��9�g�g�3������|ڥc��>�f���O���J��K� �3�Ф �G<��g����~y������s�|����s Pu��ϴ�g���s_Y�v�絉ľR�+�E��F�h�j�-��OԶ�h3��^��q|VD�����s��ۜ�v����{,�Q�1���p����&,RϫW\d΅�E^�d���;��LD*L}򓟜��yԤ�K`1�;����z�.!Z��mևN{���	C "PR��!Pm_��W�sElLZ"@wD8�������"-=����W
�T�^� �DB�ig�G��ɾ�Mܗ��?��?�jg�+�Ȫd�k�����;���R�3�#�+���s�M<�O��2%�c��3f�A�"���[�G�Q���f~�nL�ᗾ���f�����h�pck4?ad⛕f�4���V��±ߞ3��KkG�o��x߰��h&;4􇹡�{뎏N�=�sVBp�"Wk�뮛2h���e3�*C��V����t�pkC21�a��z]�r�Z������Y�&K:��	�E�$t�-�w��%��g�4!dZ���6B�2?��?X���C�6M�lV�cr���?��?l���7��G����YD�=�=9��p�'=�I�����s�."Q���o>m��2�|��6R�xj��4��~��ӟ���ܐX53B4q�9:�k^�{���d����VB��dK������*��3�)Z�&�vv�K�0G.t�~^u�aj�ӄݖmͧ;"��+�&4
�f�����q��^�"������+8e�D�V����Hr?<&2��C�MU��J��Q_;횵�Lov���I�9G�� v�/b|��V��ޞ��t��6����
=�^���1��z�0��8`���3M��D"8�ːp�gد�_;�Db����өC�E�w����ɟ,h�6s���H�tJf	J�r�]�j���U;K�gJ>�\�w�jG���(�:�Mb)Fnm3i\iZ�MEq+x�F�oƂ����u��|��R��C����=�Π�*���_U�z���j!�9�"a�y��;0�,A9w��x]�Ʋ{�Tx�|f�i�4�B��n���&��ϴ��c�� �ڎS����и��+
ә7c7�CS-���&���h$�h�UՇ�8���Y6��]��[��NmNgf�ʛ��ߜW��g	��P�	߳�9:�ϋ�!�	�~�}�N��p�}�!P��ឳ�!d��9�<���u2���
M�sʕhmV�LI�W�0��=o� �����<T� h@���f���:B2p��`QbrY�6�Q�i�L�,�I_�r{�e�i)HLڊ53d���g�`���r���§�6y�g�������l�;�<��7������ʃ5�p�#�򾦨�M�}.�5_�}s���t($� �Q��v��W�:���2Hw8����>lrw�r���� �������nj��,A��9�\���Q��ʛ%���.�!�������jXm���ѿ�g��o����x9l��`9���:�>�Ut��G�gݍ��{N��B�{�Y���i.��I;n�B�Tq_]��}�B�b��3u�^�1�Ye�� �\S;�o��1�����Jm�>��}p�f���N`ϟB.c����p�ĩ��#8���ۮX�G��_��E�m��0���Ɵ'N���:El�z��C�[�Wځ���������O�o6��@H�
(��#���^��gQ
�d�4C̚��T#s���F3��,L��U֪?����xS0�M�߬�����57�!f<�QR��]���&���|� �@�X0��(���-.�i�2t�"K���Zf�5������E?��,�̉y�y��xl�.:(�Nw���vk��lU�MlX��c���5�=(��{?�o�3�><�.`��x`,�/���åJW�g0�H�K�Q`��[����x�rY%+�O�i��N�ɬ����s-��~��2J4m4��`GmT@&�M�B�&�	�̊�j�p1�q��fۛ��\��!�+�k��7��}Ώ��E��������?��D�T�Jy���W6����y �v�)�3��1�:��@�_5�4�0�,X����J�����(�r9
�Y�9☣#���(Q��nc����u�f���$���Ex�&��oW-|j�ϴUVz�?��&4�I57S}s�s��~��e"�ݿ�w2�5g{2 >C�2LG�Fĵ��ZLG�舮j�D��h~�F������ʢ`C ���O�8y.���^N4eg��Z�ǋv��s�S�h?�<J�-��<��գ���?���������FG(|�9���Q���-K)�چY��5A�)B��gj��>Ke2�Dg ���K^��/3�Ĩi�)myQ'"lGC�	�"���U����F�������Yk%iq���-�poT�-�r���������=G�f|h���8�d�X`l^��;�SJ��=7=���f��ZAo�ۋ�&��	��-T�^�{Eo����/=�
*l�L�.{�#p� ߯��B2<�'|*�ʈ�&�Z������o.P��Ԝ�����e�b0N�������O���t�!h�P�i���<�'ٿ��d�x�[���t�ME b>��k�����k^���6�Z�֋�NJy�y@FZ�}����T�1��L�X(k�A�_�ѧ�7���T����˄�t@�2�|�䳎tqBԦBvT�cy���٪� �^�R0#����� �ڼ�v`OA1��>���
C:og06?�W�5~�}�v��?���bC����N�-�$�����P:�r¨T�m�p��۾��u�ٜ�F��o,�h�(�XC��y2����V$l�En�äE��2�H��C�d5�ְ*kB���>�<J3�Q�}`yO�^�	���-��@�@���f����@\s� �T匚�|4�v.�y�.�4M[9����7�&��O��V۝ʱ���s�����#�A �!ad�=Z-6�V5;�z�[� ��I������pТޖ����j����V���V�A�c#p�fפq]�`bׅ��i�Ө�=+M
�����h��*��I��@��G�o��h&���� kRNM@������M�]ǂ�W�����i��N2�j�Ь�DTƣZx��07�
c���|hz���}��i���f����]��a�ɲ8g�	G���?��X^�A���w|�\B�R�m�s��yF��3���:W������3�Z���w  ���,��u�ˌIx����#�mv�X���j��;=�\r�
���b�f�����l�����6����VVWoﭮ���6ۡ���������p������m��j��+��S뽕��5���i�;;��#�7 `�A2��	�l2���5&�G�T_p���*�I
��x�_}\�cQQ��X�t�+���ɿsҙ��9 :P��j�E�u�tMYD����O|b�7�aϹN^�Wۍk[�~��㢌 A00��ء�i|;�n���	������_�*~��#�_d��\� 7�P����r�"�f�X��v1R�b6�Y[3W����Dۘ��&5P�
f}]�އ�%��9��bѝ�H�`^�"��k�g��m�k'��ub����S:<q��m��S_X;ٿc��~��Be{pb�3ē����G�Νy����Sw67?�<zg�������U�Q���';E��q`Pj;Q�l)���t]A1KT����S���*t��,�嗿��͓����0|�[�ZTP.�T�W��_J��I&���,2�yf�!ϯ���'��֎Ό�p1L4g�jީ�6ե��%��Ї�Ї
o��u�+� t��c������O�g�9E�:K�G{Ws�}���'���?}"��'��yâN^��m���  G�\��d�A�ӋBY��P�m=6�����@x�I�Y���w������^�������m���W=䃽S��sW��~����}��Woͺ��7�w��ӟ�X���U���Ǐ���g�~v�̝�\��~�a�!�ع��g�_��Q�dK��yلt�#DE�:�p�Y4H{h�MoFmReco.���;<ݿ�˿\�b��>�,�js����p��F�^R��tX^"�e����?۔��*o�ڋ�~�2��~����0}I\�/��/�=E��vJ��K4~�߂��|�0��
Jx7��E�6��p�s���31Ͼ�[��h� b��)��
��=�s'�o��oO�AF�dx�qҡf1afTI�o��!����k[�'O~~p�C>�y�U�>����g7��I7��|F�י����������?_������o�>�՝�����>��1��Xg�G]�&�A�ƫ��1�9�����_}��W��`l����jm.�����8���>�,�(��o3Ѳ�/�2����p���z�긓>���x�R���ߘ�@r� �qcƯ��l���4f��� �g]5�״�BڬYl�M!���E�"�se֣ a����0��PW�Im��� ��"��	��`Yσ8�<Nx�<�茘Ҟ���<-C�O4�VV7�n���֕y��UyO�a���O���es@������z�?񾇝�����'���yp��ן}�7��5ɬ+�dҍ+�MPڴ�İ��F+Ӻ0�[Y��U���:����Jʤ�;���
�Y�9�<8XP�x�ɬ�ʻ�L8�u/�^���$����\}C��&�B���{�)��Vp���l�"{�bV`)���ؤ&/���3��50�]_d�K��e�R�y�o�PTô��8����!g�S�z�э�ŝPCR�+�^XD��1�e����>���2��S�G�	���˦�&G�.K��y���P[��h�����8��s��݃��������}��s����?�����So��/6���hV������+7��*4h���v5�W���_�����f=,��$ʢ�g�����ZA��ŋ1�:��Q��D�:��^&m$��«�C���6���Ѱ[!L�v�N��2R𤗹F���Y!j�'_���8��Ƣk{l�7Qp-��]��y����1HMH�X��6�d��BH�b%������)�B��O��O�1�
J'S�^)�f����q|�jkj3�A��f�5zh?!`�ۍ �������<K�]����C�e6`nQ ��^.�z�<c��9�6:"i4���������t�ݜ�m�������_y���C?��׿��8�������/~�CkW>���F�ίYkzW�{L�Qz;�����~��8Iz��W�cw���ʇ4ḁ��l'[����؛`2P,�N�y�BF#��UY'�s��ܢz"��&�\��
�+��d.��ȝlf��f	���RsrմL��2��3/{>��
%��k�~��R�ÏV���L����/�2 �dLX�+^���~�Ǧ��2痾���ق�O_�QD�=��y�5Ρ��,��c΢��B�9��w�wO��C.�5�����/�����i�maԻ��	���l������s-�:u⏆W�~���'��/nx���1�-?��}�i�����`�����\��5�vm�[/��j�;�bP�K,�����|Q�e�7n1L�BH�Gm�fM��h�+91����w�|�+���+���#g��.θ��L�]"��Х.d�Ѭ����P-������\HDU�%�	K�"��^\􋠂� 8ٺԾP�����7�\�ז�(��HQkk�ׄ�y���β��"a�-����x�k^S�jS�AHsJ�f@栵34��X���Q��Gl.���j�_Yk�������[}�G�u������1�����������7���w�����7�|F�>ͥCc9ܯ&�pƼZm;��xFab:�TH�1kJ��^W	[�{v6ÄX�l�|�:"s� ʁ	ͱ�`�~��KFcEO[�ahV�X~���c���}�s*���lbR�Ǽkxy��	� ��Ř�)a&~�@��)'��3Q">����j��BV�<@˃�A�%��>�N�����%�A�_���xz5D��i7f2i������훠�᱙#�Q��0Zoz�'ϵ�����?������>��+��k����:�I+۫덆'��z�qt�Q�+��F�J֞� �|�b	�1Y��v�%]�|9k������N�L`������L{��f��]:K4��%P갠K�RŮ�(tXD��<s-�<A���sSP��=Hm��P/Y����wY�s��� m2>�!�KPt�9�O�������p���f��F�)Q�O��@^KM�P66���_���1�>�~�0�ߏ��Go-�-�ڇ��F<�/����=�~ss��7���'����GW��9�[��~�~e�k�hX�hkL� յpxY=M䒔�c t�������EH'w�5��
��|
g�.*�Ӗ�m���1�����.aH�h��P����&lȖ5��:�vQ�)L��&<���}Qɩ����6�%@�
�.��������9>��@����m�s�B����z"�Ed��@ �`$�>,�98��>ۇ��h%�$�����տ�Վ��3X?�?6O�x�'������>��kk�>}�7�����`篍��2
+X�{��E{J��1q6YMlĮ=o+�&ֶ�M���%9X
\���SebtCdtr-�I2�L]�EyH��ѱ�%��`wCxX0x.P�QT����R���j�zm�?�Y%���+�.�c�V,ͺ�ـ���O�I�L� R����wO�]��귄���h��)�G�`d��،E�HF�:7Zլ���|��˽<f�7,2����}��U4e����Y�F�n����룍Sw�_����ɵ?k�c���_���'�|���A���͠z�'���kE��}�c�⢎i }� ����sY��\�A�;�
VO��vf�>�/�o�����ȝ!pȩ*v���\��Q�}XA</�������2+�������&������"�1%���a��ʐ.$D�5Gl�'�$�߬{��?&�5�a�8�ۺ
A`E3�&!��I�hl��qaX��25�,�!�b�@x��n;�����`XP01^�G��&t�q�c���� ������\u��'�z�؂��7���a}�����m��k�VUMV��N769�C$���K���-T���:Hǂ81�����b���$�)�c�Q�Ҹ��yWgse�a�ߨ�˖1u��lzk���IO�hٰ�>�$Fp{\?�2�5�@�'Nxۤ����!?NJ�������ctpZ�ŅqY���^��F0�k8�ue�H�X��E��'�s1,cK袻m��rA�]D����������_�k��5�3]Y7��a�f��7h@�]�ɺ�j���?������X�MVȲx"��{��8������Bxp�Lo��.�������k����$e��++��N�E��~oog��a�h0��������V ����1eƆ�X�(D�M[��ݔS-�z7[B�s3�;2�B��Y���jS���߳��]��\ՙ��q h�:�U;v5Na�=�+�<�XQ���gϻT���?�JAg�%��u��l4H��E�3^,���-��@ծJ;�����,���R܉�Y�0� )���h<n��ŋD�P:ʠ�B��VމYw�E���pXPh'Z  �hX���C�7{�:�4"�D� X���w�I����I��^�J�������-�l�ߺu����DgO��w�ε�{��{)]��:��	1��`�"��&Ӹ����)@a>L
xuq,�P��}3�����L�aT�5�!�,���.����H��:׈̐&"�ﮓ:��tI���sml�81��=�=��y�ѥ �]XV>+�8�9r1�8XȌ�YV���׾p6��q�Oe���-�9��|D'���G>򑢲c�!˫�[A�+���H[Ԋ�%����E��FD<^�f���C�-`Ig�<^��M���nIu�<����\�?4��W�7����^�k.�nN�������B�e�$S�����%h۽1v�3X�����3 Z<��Lm}���3S�r��tҩ���`�d���U�d����@�.��䟌Օ�k>�o*��%�f����T2�jDs)�Y�M�x��������3ĩZW`�"�w�g
/� 3�Q�[�����E`cG~ӛ�T�0�������8�>�M�k�4���j.�>�s��\҃y������C�����u�ڡ�f�����Ͳ��C�{2wj'�QDAkG���W�K��Ѯ��;m�Μ���x�7�AU
�*Lt�9b���d�����ΰ (�h���  �3�|��nGt�(��1�Đ�b��,�D�n�.Ѽ��i�E�h�캚�!9FX��\���\��k���)�J�J)�ٯ<��3jf���������N;���#2US��A��A�8;3B��R��{�w��r���cN^�9�ݐ4CE�.X.4���_�Q
�@�w�K{��q_�s�>H��:s�r�>����oIZB'}���]�Z��8o�oj�mtP^����6gϟk�7w��u��n���X�q!WhQ�L�<�o��Ewjǈ��w��3%�8��f��	nXS^6������4mc��ն��K���ڜD����J��մ��E��T�Q�=��nl�p��U��1�Y��EW��w^�WcsQ,�����k�(��.�FZ��h	(Ζ,Ma\/j�0�9#E���]n���U)����0�n%Ys�*0���67�5����Q��.vd�?�wv'�`�[K��Ɖ�ϱQgF(�\�Ex2�B��PX�nD�N�L<Q���N���zO/z�	���qMuZ�bׂ�5�3��U�\�ḿ�lӌq)�$jS�@��*3~T!�y�ť��86
�T�6@`q=�-�s!y����F�i�{-{�qHZ~Ja�(�d\\d2�85A�a�^�v�<94�qmHm�y�}LܨX�;}<s]��vv���/e�;� �V;�KK��8��Op)�n�C��B2İ�ӻ��n_��t�Wl�ﾲ]OW}��h��zŚ��u�9yb\����얦��k���6�O����Y�r�2�,y��X�tR>�Ne�I�3M��5�)@Rșƪ�
bJ��bemUX�>�̉���&����'�Œ1�
)��M6A�]�KCyF���(o�;�S�)L�\8���9j�>1d�J���|�}��rGp�s��!�O�N?F��8�|��WM=���!&��7�����"�;�`�~��߅�-��Rk�2I|hW��N�-K5�щ���ک՝��lJ!��}u�l�b��=o�����iVڱ�z��f�?.a9n7�_h�����y�U�ze���kǵ%B͑���~��D
�Q��r3BU.��W�WK:�ꠅ��頼_M5�f��~��|�Y�����ɘ0�uT<�H8mԗ2�N��3����i����C�{�!f)D�Eϩ~f�L��-o{�ۚ�����X򥱻����L��@�E�<pw�)of?)�r;yy-#0܆`f?��8=���:��ej�fa��h$�
ND�vk�Ȥ�Y�&ΏI�(uo9��N�ܐ1���՝�W�v6�����W}�E��}L�;mek�-nX'U�K_�vƥ�餭���1�	��i����|3l�J�vONd�	��L[����)%ӊ:-��w�I�'[U�+��Y"0e�E�:Lތ���)��>�L�^tE�])�:�uĀ�a3hG�8�$`{��ҟ�fι!���󬝒�D���~5H�l,zj^�gTK���"&�s׵�Y��t��4��?5O���Y�n۴�-+eN^��n�������9������P<���7޸2��?bo�����G�b8��XN�Tk�V+�W��ca<)�Xl`-���L�� �T�e�E6[3������L�a�rɕ�Fl���TSiY|kR�	�ʐ5ⵄ⥎��t�9!y��+��LB��/��4e9~VJ#L��<��$�m�1m����?���~�2�NH���z}ۇ�i�S"���t��Z�,���0��d�q�K��~����9�1�_γ@�7��	�T_�.�M���y�c�C��o϶�̭O��x�Sox�g�n��G��[n{�`�oX��z��p��S �v��={g0*q#'Z����l6'N��
K:[���n���&		&�� ��E,��'g�&�B�(�(��oJ�0Y��qN��6[���ښ��7(٢.��3.)���:4���������^"�4}1$< ��A#���Fiy����B�*�3�7#���1P�1�����W_����d�l�u�!A�fO���:�Ut-�ʵ��_}�u��a(�Qɳ9ޔpg�:V�(hA/�:n�Ȋc�z�L��k��Z���湝ǯ�{�3������o?��t�����k[i�5+��IWK{�������q����x[txr�9��hΞۜ&R����|`�	�gr�s�A|�63�3@���|O��QM�U�Yq���t���`ڃ���q�v����Xe.�
$���}�R%�!ǖ�s\ja�3[����a��?�X�чSM�EC�|='ۚ��4w�	2"Pڥ=^���w��S�UѪ܍E��-}������ c(�ǟ�n�s��/#���ģ^q�"vX�E,�cBA���KKZ�K��^��8�4�L���7��S����{�I��g����n�����ǭ=�Qͭ�]��u�	+Ý+Vʆ�Â�K�{ㆮ��0��j�`�!���:�ew��1��wu��g�&���2�67�p<dc��Y���r�6+����</�-���٢{��D���y�g���R� ү�ў�����1���@�2ce�~A�6\ZO�Y%b�����{ɧ.�6X��s���cjU9?D�"�j�P+�gN���A$��G�8�wT~�\��Txjrr���>�*j��'{�������Qq�x/K8�joxf��;�y����x{ȁ���D7޸r��_����OY�����!��m����R-Z��C���v�J��F���V�����g>5a�a����0�^��WM�����R.7�j9����ľT�&��ZV�ʭnCi�K��3�A�@��0���,�d�/��,��Җ�,��)��Dڼ3\K�flo��B�q *�%���X�y^�6�ϐ*��M���وP�
CFBh�b7g�0��n��E�Ĝ܇ҕ��sσI�~ꧦ��9A�u&�9/2[�=�m����<ƉyTk
a��}'ьs�����rG��h6Z9vb��Ki� ��Qg8h6Z49��z��]�|ss��w>����^ks�
�}⎧������{�z����ںN�I4�8ך���Ѷg�}��hՉ�v�yc!Dm����)�Rq�\}3��>�^�Bȩ��(Ԋ56��`&���ht�Π���&`V��v>m��q- D��/�lE��_L�h��?j;fF)ty�DN^���A���O��6�'��6��ΩN���H�
��d�M�cY(E�)K����v$1�!\��S ɬQ�T�KH�����nsDQ{�0�uY�uu)`�&�v1�0&V6tN��c�X�O�*��Ѱ���ޠ���������i;u�
�a����gn���S�������7��?>���Z|ݟ~�/����/����x����+(K�&��+po�LG���]��v��y�7壘�D6�3�©�����Pb5k��P*�#/��mͲ���|�̧J)��ȳRHUJ�q��j;�1�-C�,C�	��6�@��E����h��{�Yז��ꈊzLs��̞T���3�*I�1Ρ���uf��c��9W�N����]�]���z׻�Ü���ٮ\�R����	�r�1��t�M�(�u��i�����4j������[]+[����Q;N����͗��h�;9>l��۞������������w����O5G@W��3'N����in��[7��E�v�>����:��~ �����}�mF�gt�T��.�<�Χ?��� TO:�dl(F]T�ļ٤k���0��&`��L~��ɉ�3&��E$'oz��=���p.��E�BB�f9&GL,�:*C�xT&��M��qн��on^��וJr�%���X2Ь?�׹�V���o"<#�����|Ԙ��Z�?�ݖ{���aoeg�26�kK�o�� ���ŃV�g�;E4���#���z�+v��!?�Ʒ�x���=D��k~�M������o���7����ۛW���ۓ@�X�܈�"vx������͸��|�T��F�ZO��R@�z�]�ݵ���|f	���11E�:���oR��!Q�IJ��	�|�/��5�����늶1�Y�1��yη�LEN�./Q�6����}���0��~N�0��-oi��ۿ�b��pNa��w��1�sc>!��(J�v:��6y���< ���
��;->?�vJ��x�L2ϲ1�p����J�P�w{p��w>{s{�����#����_{������������s��So�q�\󹫯��/Y��5w���[�~j�mQ{|����~��/���wƏiGU����Q��\1]���{�ʉb�if�V�J-"m�NLQ����N�����$���[Ln�M|���,^��j֤�oC�f	�㶩gy��\h�q��(�4 �%�[�N܃����#?�=���ȏ�HI�f_<l�V�s�K�dF�8�� �9����.��L��j���7鷝�س���6	�\�l�����R�E��e���(��IY�5��Xȭ�H���P���Z�w�k�޻}EsŽ�w�=����W���˝��w��_���w����o�f�8�~�n����qjcutzx���z���YW�u�3N�{���g�y�����~����vo��=��`���a��P� .	��������6ᬠ� -S�t�
+
ΐ��E�t��愫�&\n|(�y�Wz��&�	�S)��s쑊�&C!�4작���A@3��]��k�p.b���&RDș�,E;y�k����YD_�a��������[+��	�Bg�a:��o��X�|����Ú��,�T�ﶝ�{W#�Q����gvg=럍mV��b#C�#%Ĺ���-nV�H(\r@"6HH�K�,$�	�A � !���(��8��z�;?�U�{U�zjz{v����'��������W��{Մ�q��ѣ���EO��VU�*ݒ\<�[Q@X\۵+���0CceB�W�3$I��Fl�ɭ���R��^>*gO$���hddf�HrE�M.~�o��^�i[�Z�<���e�I����C�4;�,5�'���Q���PF���=�1.h�%�F������zh����XK"&t�@"/���m�_А��2�]Q}�MQGD�D���K/��E�W�ԡI���|$ȓ���(�>}:'�li	+l����Z#	�ॲ������Y,��PG�:]J��K�U�����}��j�zA�H��G����9�`�$�'P">t�P�lI��,(ݢ�IS�lH��Z�u%�S�oBu������ f=[ȹ�S�/|���$���ρ4�'��0f`�`R�TSHÅL�D�Jq����+6� A��D5����cB`�I�U+sY��(�y
ucB��\g�h$u� �WR��P?*�a�@�u��4;��9�� C$	3C��^;���`�Z%��P��,������/�B�Ӊ�}�a�t�~�!_��gb�'$�F3>DqUg��_��A�����&w|����'o"�$9�h�$LsT_Ɂ%D$�^z]�*��"��(Ġ��_v�����Q�#�:}#$e,[tLB{}�b��%�*IȾ�M������E�/LH��.\ )�����bJ2�?n&ѿ�8y<N�Z�
FNC[5-������a(u��E���8��x�ep�U_D�i(�Lڭh7Ƞ�3&l��ք�d�����R�cf�"�����+�2�5;���J���\]F�垅��sd��}�Z�_�����>Ń%�$�~�,|H���r#h#m�&�N��0�=�a��!,w;$5�ݭ6�+vOKܓZ�:$�:zx=P�g%�Ǘ�}&�!����Ɨ:'�Dj؝4���Ȉ$A$Q�u�e��qHڤ�݈o�l���y�}Q�j���^)�|1P�on���߈�I�e�쓳��`t����Ե���$,���|���b���Z��w[O@��Z�yh�PYG�*k5qKP՜%7�&�/�<=l$L f�����%�Ђ���V��q�q�Pd��R�}x��5/H�x��$2�8k��*'����q�U�4v��đ�L7�V$0r��-$�����m�{�( �M5�����L
 M��TK����#�@�
LIe&h�բ(1^�ܶ����F`5;ٮw���}�Ң]�o��ە�k�B���ۤmc�7�� A��oޯG�_~~�?��'�~�����I��\��]�>Eg�S����Aq�A6��<B�R�����?�䓿y��W�R�UIU���O>��w~�R9�Jh4��.JH�>[�\A2t��Z����1�u�"�J�
͜K4��ƨ{�&p��S��њ{i�Φ�i�X��y��u�S6��T��>�|n���k��Xa������_-5��
�@�;���{(�=��r�F+�(6�.L��t|��͕�F�ïK(�I̋1���l��� ᓄOt�ٞn&zIz��z�[��F���|�z��I�4"�dgMs���o=����:���b<~c���v�>�0/���]��X�F��z��'2�2�vY�ב�2�% �,y��ƥ��:�.��y��2��WweŘ����M�Zv~�4e�KR�pz�!cf�f#0���s$L�������Ҷ���TM�r��)aI9S���U��(�߉9�7�@��E+�L���O�E��v��(kk������ҍ^D�Ϟ��Mb��r��e:ύ�|W�2K�A���H��<�*�&���bؿ
D�H��x�g���$���^�9�ƛ���H;m�MYzTe|�F(����d̝����a�bFf���ˉ¦҉��L��W"����N�)Cʖ�P�v)뤬���|�����+��|��׼������n�%�N���&Ν�;/B��N�|?љ�T��0c�����D����̩+� ����H��fLnI��&�Z�� (кo2� a����:�A������,�{���ܢ�����?>��S����떂}�������?|��Q�[z>N���1�b{�*5�!s2��*"R)j�'��b�~��v�Lc]���c���-�9q��'evQ;�w�~��V�LsI��/�'�hێ:��V �$cn:͊v_IG�<���V��� ww��(k$�A����3�aK������0Q�D7C=�τw���|��=�Û	mgV�/H)�LLL�=r��/���9v��ۈ�Bv�ң��S"b��hvi~�j�>[��x��1Wh"2C^��mA��r�1j�ʎs;�k�QG�H�K���F#�褶p�ɮ8�J^H֙�S�Ga��J������LKnE�|�2f�%�F$(�k;�e�ۦ��u��J��󗤺��-��k��i�Ӽ��n,ȵ�����p��E(�k�����b���;�Y�!`#��>�j v��|8ۯ��Q&�o$��h�Qy�x+"7ȹ���Q�V�-�7���ܾ}��<v��^x�O6���[�OO+��'��F-�}�+s_�K��h7�<"d<�2U�*�@sM7\(�y%�:�� �I��u��I�ܑq���KA�+!gn�������a�0k܆�]L�2W�Z/��Z9�K[F�Y� ʮGm��	[� 8|]e��i:�U}�ݟ��M���r���3�C|��Q�r�5�g:�	�`^DѲ��(��qeTF��
ɭ����$���x��M�<@�ve���o�t	ig�.�Yv����B�le/珅�k{֑Վ�g^q�U,4���E�:W\_��5�z��}tٟ�A��Y�.��o��Q���j�\~�#���FGG[��M��?}�����O�����_߿�={���=�3]x�[7��g�V}��lt����X��iV������{Դԉ�d�ⱝòt����p�t�)T1PqUe��E.�a�P�]>�9]h��k�/����IRvS�	\�)��C	Fl4��}���FSm��n�.5,����r v��͐�� �1-@�7����/
	�Ur%��@q���r!��mvg�င���+���(p\d�G"�*V<�Q4�rҍ8m����92r�Y9��t<����y�N�8�nvS;�l]�#|����,;?x�F�V�یu�a�y���=����x	ҫ�j��c�=V�8r !G%�T$�2���E\D:DR�}^�х��l��,�����7H�������;S>*��r�A�%��|W�D����D��D�8�@����^x�"�v�DĘW�	Mb@�}�����d���Í�{n�̙3l��>�R���f�:���7>UK㥆N�D'�v3*V:IAք&E��ɉ�<�D�I�0�x9j�Q��	���$uǪ�y�J����ߝ9>=���٩)�N�T��s��_a��W���T~�����ۋ���v��N��u��g�u���Y�_��SǻuuvV�LN�=V�KH��5���|���LMIv�<:=][����L��Z;Sz)br9fzeX�>���
i�d/٘�Sc�gV�G��2�>g�k$�s�ߥ\Xے�8M!���Gؿh;� a?�}��ӄNT���+�J�b8�D������_����x��x��ָ�����C�ML�����Ǒ,�-c��Eh7@�}�СCOMM̓���AE��y7HV��z��M
RfN��Q�^�a���9�_fl�������M�k6��l�������~���͙����by�w�N�=i٨2]��S�ɖ��,�-���I��2�!&3���]#��X�ZjT�� ���Qm��e5��"������A�w�n���V�&z?������20��(����k�g��Z���R%�@����Oq�ʝ8��@r���
�U����0^,I_(��r6 �
��Iv�����;w�Lϟ?��8q������4<��U���v�h6Z���.^�����{wף�0ȵ�H�E%��@0�SβD#Y%ZF�8 	��L'@2F���r�w�Q���Z����DfQǑ�*"IϦ�OQT�<C:��O
�Y����R)k'i�J�T"ɡd�h4�������������{�l	oA=s����W���.�-����إ��y%޶��l~����6ν��<y�d>�1	�t�Az�F �-�	V?�kl�0ξue���NS���N׽�� �7`+ ���V��V�]�q������e�!k ����v��Į�I�ㅙ[���/�����!��������GD��F���w���p0�UL��:�;I���ή
׶/r�'��ga�dgaa�llafbbj�p8�R��hN��҄��


	*2.,B|J�?���m�X0g�?x����sJh PK   O��Xs!��}  {�  /   images/330d02b8-4530-4fd4-b6ae-26fc03cafecf.png�g\SY�>�cAQ��� *"�Q�Q�t�ё"�"B��HG�N���'�(�.%DB�HhI !�?fFt�y������0�!᜽�^�Z�j{�]������^�n�����[�%�n���-��ߘ��I��z�73�u�,/����:��n�Ⱥ��Ս|'zJM�~�K���?t_F�a�ŝ6��<�x������ޡKw�Y����֡�i��WOt��O��3uF�.�?Jh;�@>Y��_�#�5?A��ۙ䖥�R�L9ɞ�*�4�?��Y���ﾫ��o��Wm¥nL�n�k�R[�a���u?�qxS��ҝ����RR�T�"�n�����oFio���?�q�٨�S������ׯS?���Ư�[��Е?�)QAcek��h�o&��쏮yAH���;_ߙ��N7!ѹ�/�m�߻�����3�ֈB٘�<��%�j�7f }�KZ
~~,ۣ��ˋ)ybz������N� �e��A'���ˣ��.oH���f���ʞ4xd$�U�<�o�z�1���ڵwS�9a����8z���J�2���y�u�o�Pyz`� ��b��*o�G�D۳��/ep�cҘ�ܮ�%=W
��c��T��,s��;���#��S�'�4��,�)���\�jR�zK%�p+��5�'x���U��u�G�Z#����>���ԇ
^�x�6<H{��v����"�䫇�Ed��U�+'B��"�����3���O�7�65�_��E����1nZ-Z���Uލq�Nm�ě�}�̦�Q9ec\�PsV����퀴^��>l6߿ӦИG3��	�BĘ�����p�����v	��I�Q0غ���6i/Y��&��7��vJ��x\��٭2z}�v��H�?nP�[�#�-�(�'�=z��z&�l6�xh����/�� u.�d��8'��H��/��m�j{���$�E��M��w��A�7��~[���IФO�-w��$�6�^�!<�l~tyu'�i�coB~b��X1��["�c,C��ň1s��x����3�󽿵*�����G,�7]h�4��f��T� m)KA���~&��G�g���U?�����ų[�;m�|�DF��gS�dD��Ŧ<F9E�d��ݢ���J�����홈:y�U�fz4�&���ھ7T��L�1�C�����~�����K���q迪�_�����6��!�H����4+<���F���֢���7��ߪ�)�Ѫ�dSW�.��<��[ ��)�/��;D�[�Yfŏ%}�z���K��:����m��q헊;�����>P�/U�C&<d��]=�!��1wڂR����-�J��Q�r�>d��E6P:�L��^Mu~?�/�|X}�k�'��6ɑ������]��hC_�����o�	�.+ae���v"m[m����5muk���}&�n=bx�c��l�	αck�~R��'��ǇB�G�������1���R�`�_X!8��7�v>̩U�[.�8r=Uz����ȳ�(���Ll
���<�IKj�~L�{vl��|<�k��E"Vcɳߦ������Z�-.���m����k�#S2ڃj� ��ئq��9����6L`۝��/7�͞L��(�0 �R}0�|0�yX<����G��I͕�v�?�Fr�����t�H^�_qLt��{�;]v�q���1"��	N�����=���������1��ú�7;�ffE΀��`�������B�ٻ�1�D�[�kx�:#��� j�/�:/}���PR�c��t� <D`��5�H슛V4_K�������e���0�#mu����Aڼ�	E�H�a�����7������-2ծ�H�?FU�{���
+˹q�ѕ#2���~L���<�S͏����+ �q���?:``�',�:�����{{�Į8!��܏�� �iC���\���©x�//�h_�Twj|�`C����L��OD}^m�z��i+z�z�P���l
���0g���\��Pw#�x�E\> ��E���]qGd�V�=P��+��:�ds�x�䷈1;j`؏�����O/o�����׺Eॶ|t�C��i��ZB E6{�z����πsQ<�C�;��䐘�V��x�����]����g�ͅ�M�iB���=���Pƥ�C��T���B������D�=�=��I~����:���19v� �;��~tL�o��'���B��!Y�k�c�5��WZ�D��f�܇�^^���8�a����YB�b��'�"�?z�s���P!^�IRS��p�t���6�����=g�C��k �`�A���|��%K�����W�����U��*���
�_������>�'��>��"HO�8���}J)��ۗS>���d�]Pv��wl©+���qݓB��zj����:J��$��	��pwQ	�J��S��0B���w���І�-��(.uBſv���"k��=8b��IPZ��s.��m��Z��iyb[b���fޟ2�]#Ž��!�}=D��F���<%D%��Z�xڼ<B���͒�>J똵�����q�ź��e!��ʺ̘�!�o�%��h��9��l]J�������|�"�U�c�\0�D�=�z���&f�a�唖��F#u�eNY@�Mc��~$'z
i| �k�w�Na܁{�1�c���8�r�)>.޽�kcN6���ʡ�wh�_$uL`�����Ylhય��J��X&M
T�,�.�1��־v��}����^�|�B~ν���3|�]KҦ��2�G��n"a�QY��е�G��Ӱ��'D*%�^<KF`}>�]�F^� Ŷ�1��"E��p�K�Ot��A�B֙Z�������a�w����r��\���8��Z����Qd���(_7�/$ת�f�����jQ���D�2ݨ����E-������)Y^Uۙ�B��nٽ�^�Ǌ�pM�H�gG!��5����O�9j������&���·,"�ӕ�j�w��4��z��kGSez����]�X�̠3�I��l��<��W�o��s��!CQSx��Y(������rw��ˬh\E5��Wt��̓��9k0��d _��ײ-Q���xfr.2��/8�� �<����G��?���]�9f��S�-E������6�Z���/���ʶ���h F�(}D&iKpi�g��??Y+������X ����v���s�ٴP��"�ϥ��o?�`/7�l?~�oJM�=b�霤]C��Zu�c��@Wl�B�~d��Ԗ�¿��Kk����F�����h `VХ��gL븖1��:	X{$��6}"���![}��#h��LŎ��#̞�Kk0��?V�=m� ٥�����o^x��I{ǈ̆3TV�����ŏ�Tz �b�iZ)����<��#��\�]sn�/�`K���2�sq�f9��)�+,�c���F^�Q5�=e��!-�[���q2�f�����g}�Pr�)���Lj]H"�л��隶��Yl9�J�����kj��>����Gr�zGg;B?������-�{ײ�3#2S�$h��d�Y[d�<�/+��qԹ��<��Ι��T�O��ħ���ලl�~֕�6KD�}��.����H����Ԭ��w
������e���ǸÛ� ��؉�1���{��pj���{����9���>L���O�8�s�1�)�_% J�R&+�����D�M���þ=��\"+~���Q�r}�Q�v��f�L�e8��:Ǯp�뉟����f��>���c
5N��p�4u%�n(B\�}��g/@:Q�h�`�piu_g�q輡����婬�?*���gG0kx��?�����s{��_�n^�L5t��6�G�N%,ؚ'tr�Ҟ��S=b���@��1��(����F����6(Vc����Y	���F;j��Q�'/T���Dv+yA�v��}^Q�Ӹ\̓�2�)g�\������&�w�����a�1���i�l�ZKA�S�Ez}H��D�,�Hr�W�}O�E2�R�R!W�X:Sm�W^^���N�d|%?�W�S;��*;�Ayt���T�u_eI;�><7P����ɶ�E8��E�iఙ�a��I�D���<~�Į,=�$�p]�=	7�H<�G�5� /^��[Q�u!,�>~�*nљhΜ����{Ո�nz@��s������W�{���GO��H�f.�������G��P�����^j��NA��N)��X�VV4���>U�gf%g���Λ��4t8:s��?�p����c	$�9��6��5t�䰶m&i���^�����i��.��4b��z�P��
���/Hrx��l_�1�\hoEu�t���+5��yh�8ﮖOj䦠�~��ݮM���Ġ�4�8���-���ړV�QPa��L�[�tC'	#K]8�����a9�؟������ج��f�/<X�E��ZbЎ�א)P���1z��9��7"b3��~�?���~��O�)�	3����dØ|RKO顊ThU��kc��=ϊ�e7����8����Ɏ�-�N^V�2Q$�cʕ���w|؇7��*���+��.J�k"<�nDo>�=�Xf�ȟ���g�5�߫�����L��|%���}���D���]���LǓ�P��+�}c�h�ư_l2]O�� �jH�/��y���/u���`r�it,�5�=�`o��
텳x!�[KT�}L`��9�F����f��ڳ������C�/��r��F�#�e��Ļ�w�ڼW�^�'}A~�Qp�=ͩ��U��s��\�����5Qv�����,R�	�2���J�jp���8SLEk ��L��N��k:G����G;��#a;S4�j=Mlw�tﵶ"�MX�=����)�Z�u�a�E��"�`��f��ڵ�EM�#�$�S >p�����)�b�X�-l���^h����q���| �Û��v�&U��(���
�c�h�}��.��`�G�D��d�R��H�l���y��D�����"{�3g!8�YЦYH^��Z��6Jn��>��9��:6��Ά��0"��,�g�bה_om��蔞z({q�U|�\y��n(��P.��m�C�iΦ�Ѿ����$���}�v�{������9��؞T�b�01b��W��N�H�@���B�=Lݩ�����c��I������U�_w'�%7�X ʛ[+|��,SQM&t�/���/��:��>H|�YMҺZz=L�7�fU���
�_�xE�@�<�՗�Hs@�r�)O���/�rq%��*���n�o:�K�����(��W	�J@I��v�:�[*�V��󙈮%�����;��F2����Wo��$Z��B�~�ҵ��NT�h�S��}���#��(��8�dc�T�_�bئ����4A��$�Xs@�Z��/�&�����e��[)0��0��W1��D��[6�:L���s	�ӊNw�;��� ���r�^�%{�Ȃ��]f☷�/��e}�㺯�{�bR��B�J�p�n�;������U��, �ژm��1�a��ܛB��!��UU���e¸�Z�]�����粧��,HV*�$��e�y�6a&?�1�>�?�N�g.�q:�P c�ѕB�p���B�z=�6�6;r��x5"BpB���⏚��>?55�Y���K�i�aL��CK��f�l��b3�|$��D/��g���  p.�U-��.���E��e0u%T�f#�y�����3���)�V���?%�xHۦةL��t �,Qէh��6p����}���i��@�O�01��>fn��r�vCI���lرs�!���t�[7�aJELє�p[��W��u��8[� �Vy�ի�ln�}�����L�^�2����+^��Tăx�R$�r��
/Ȍ�.���� �ɵ�A5NΘ��9�Q�����Z?�ż����+_�7Z�z�=��`'Ϫ�;�Y�%�K_�yV8Z��F���̳�G:؅Ӳ�聈,��G��φ�g�M�����ox\br+�U 9i*r�-�J{�Xt�_�#��F�Ю�e�kN��,�3�{
2?�4�gIp����]~I��&莑�IK �0p�;Bi�kP��=�[E������w�b��^�~��������VS�'�}�) �_�J�t`�"�[1�9rk7�В�P%[MZZR�T��4��yL���<�Fl����k�������va�鈥*��;т�~G~.��D��u�wK�l��R�b��8�a��������\[m |�֛>o���� `!��S�j;�K���i�<�m)��T �����.��g�ʡk
�zx"�`Z��ߗ>Je�+�0�r�H��)Ma�_��2/��#��c$y��^ݟ�zc�n��8��hKó�"�FN�8���o�$�/�, S*]̨H�l'}��GO�]4rh���<�M�����K�,ܥ�=���n9Db%59�4�F���F,s1����Z��#�L�����!f�<`ʷu�����tPcR�Jg���j,����DV���#�{�B'r��0�n+���%��Ⴒp��r8$Ɠ�ĩF\�cE�-����J���ګW�ty;7��3�:f�2I`�N_�]Wz�vH�p�	j$']���>@X�Ufy���3�C���$�B�	��'zjmI3��
}�a<c�q�;�[CܻC��ͣ��]eD���l��&oUR�=������W{�64��T�ڳU���/MЖ/q�rʁ��R2��0|�h@DD�g`�����F[{�����|t���ő�
4?i�b� ���?K�F�ik2�ُV���^�'�ـ�v��[e	Ω�����O������^ L���2�5⍱�^�O�Ea�*7Q��i���v2����H�I����>�!R��a��87��1��$!�gѸ
e�-*]���q"Z	�^�	ā�1kɁ��f�y��8pi��S�aZ����q���|�fRC�k��
��I�˜@NWD�l��Fq- ���af�}g�(�؝��á�U���S gk���J	`ߌ8l�N�����{1p�n���B���e7�h �]�����Ad7=�<V��)���Mpa�}�Y���E@ �	�,�@G��J=�S.�,�~����<��4U�J#a��o��_sF>V�4l�f�^�PW7��"�R���F3Ր�(Ȣ;�sk�ҌS��7`q|g3/���������T���#)�||��}hޓ���*��� �rw"��J|��et@��aM�p	+��U̚���e�gz؏����y�1Σ�&k�+n���WP��l������y�~�VtG\��⤱6�� ��˕���a�{)fzT�_�y�£-�]���6X�r�ܭ9Ie {r�jP@_�@%[�r�?��_½h����%�yE�;o�\��S�|�F�.k$o�qd:�$����~���µ��y>�A�o��(d��(��ئ���6�୼Hc޹[7�I+��rr!�.��ҋ�˱ϸ�S	�m�(���1%u�5�W���q��Z_[Т�Ze��Aw�jir���1g?���9�B5n�l�~�X`��?
er�q�wLME__l�*�7%�b�7��)J��bl������K(�t4���o�����vq�vqX��aa�:Z�)��%�LP��a@�]���	�����hB1jq�K�X?�+#;r�b���t�-�fQ����neP~���%���L�����6O���+�Z���M����4��,H�D�D�LJ��`��V�~u��!��o
vF����*0~3�5P*�]����f�o�x����,�UZ�>=ųO��F���~b꥜^¦GwNΞl�&�8��Cf���x/|�~v�n5�㎿h�`&���'��`�t�ί�i Mej,�^..)Q@YgW�V��]�w�о���ŏ,�!��&��L������,x��� �G��0�`��(�ab���=#��6���J}c�dL\'�2i�u�!��c�L�4���.�"��':cf�u�=��ϕ��o5���Rh�o{5�"��*\���d���?U����#{.�Z�%<�4���S���㚰�~;�L,�c'�U�����Hϊ�DC��T�O���K����U�7�UM��ޠ$J����M䊗AoV:h"��U "��)�C��
�=)�i�봖����,t��o/[`��#{����\V�")�ޡ��{Ǟ��`��������~%9�x߸ޫ�ˢ�l��K폡��MpH�q���Ucԝ��S�`�z�]���k�b���di�My���e�5����+��£	��w�asw��[LP
�K�6�~���F��b
?I��r}n������B6;��J9�bEf�������u�'DVy��ug��"miT��ׁ�zX<�)^֬! �X�
���,xyV��b1���*9�l�\Sm����)7���6{��a��X��E]��Yhy�kZ��f&��
�Vz�3����*# O�뜈��]S�|v�t@#�d�1ɧ�SL��GT��ޕGQ� ^}��p�P�T�tF��UJi*�9�>�W4��GYȵ���ä��߳��-�+���fq�}|;s�Bh0	
+ǰ~�\����5⒕G�{&`M�O�����@V�@� �J8aq�q>"wc�+�>f��������/-8�)�F�Zgv�O��X�BT�0'5t�~ڸY�"�'��d�/
JS�;I��a�z6�C�fW8F���w*��t�r�a�'!U�"��}��� �4�t����X'�~��k!��P���u�ݛ�n��w�~4]����H�<>� ���r�LEl�P�79tF��>���L�!�G�)
�*f�G������k��?x�QtF���T����0Zgp�!���Z�O*gG���)yD�=_�\�(�nϺ�&�'˞�=Q9�W`#�N�z���w���qF�ܡY�R�yٗ�A���Ox��W&����_��Z��@��I�'3e㬔)���N���)�PGƜ5���i|��EU�f�2ӶZ���sVm�O�lFZĹ|]����%D�͙i�XM�wI�D�	
����F�YqV2���3~7���^�����;�y<�F�ZF�k�7�����p�e�Ȃ���������F��0�5���$�}y�>z��k��c�P��%Gl�+�&㛄�e���x��Ҁ/��;�VX07Y?w�S?jfzb��$�*�)���
�|�M+��Q�xg�S�,�c����X����>Kk��nν^����t��1��р��  ߘ6�<��#H]y����^���o�o��f���Ǟ����)��W�F�2\aK����+yJ���>�P�GF�ރ��玲�an.=Y��2�z3�{t�Hj.�\�=� �N�M3ܡ=[ �>�� �B}���3���;�2/�)2}����.ħ�Ə��f>� 61��]���>�|0#�;����F���fB|Z��D
�a����7����͡�����0m�bSZ ���ޱV	S�d����I���&E6�VH�}U`�i4|�V��8۱?�����h)]��.�s�+�����o�/&��K��by�Y�T�>ώ��h�B����ȥ��K~z�ϣ��k��p��6�� �����PAzˮ�0��N*�ȁY�ӣNiG/�]���y��yX����e�Ǝ+	�f(�*{�Ί�;[VQK�:�����N/.*����G����$Q����;�����y�<�Y(�&"9^%d��C��C0'�-:;�f�ڬ�]��;U�E4A5���6����V�)�P�pvwٓ�YC#��p;VU��S������`3NO���~�sFl��F+���N�ڲ��*��E̜g3��6��彌C/%�� �	_���0К�8f;^���,���� �H�]�z�ݮ>�җ�s�=Q��!=�A�WC�brN��D'�9�Q��ֵU�wZzJ�>c��F�B�T?�����0�����2d^r���uV��b���� �1e�k�>���hPL��_өݔ��+�%ͣ_�t�r��dy~c�P��܊���=��WE�x�l�]7��h���>\Q����v�d�x�k�`Ul���l�ә�0�t�Aͅu�v��:L�R�^\"�;O�H<�/��~ܚm��l���o#�~LF��=��6��|��\US���]�f ���ol�埰-Ev��V�6&�3p���� ^�*�I��<i��~�0�Ӆ@�մ4�S���t�tY�FƆ	i�B9j�p�]�}�{�`3:-4�ҥ�w:��FR��jP�.���(�<�J\���
�˴��J4t��gM��>���ԗF6SN��'�s=j|��r�c��V��� y�#�~*�;h�$B���a"+�F�C�9��lE�$�Ai�ǣ��@�"1]�J&=�r���J���ս�������g5`W �&%q����ץd/�ũǹ/%pZ���pI���*C�~��Osď��^n@l/Fte��a*�pl��x��fG�S���	�>%�nZ���E���Ҁ^7\�ǖ�e���=-�~i���4��!R����6I�R/!=M�r�xl�W���#�S6�6��D(���������/f�S�.���1'b-�R��}���ޔ��긖�3��$ ��z�K�JU�K$�Z�Θ��7\ZR,�Ν��C?�^�sc��&ˊ�_ɲn�U�K�G<
�;�
U_]��Dd�hY�/��<����^�~��M+kd9�ն�*��i�ͭ-+�z�E���"��so��S�9^�b{Չ!�܁�p��{����i���Bݵ�X��,��3E�V��������?
)���d��*ٟ��?��p�{���=E�	2��'fL�$j��=�)3�����6q�xWV�������Xj�vW�*"��dig�J�ς�T��fj!��ҏ!�S8�7m�n��jXZl�g���k҈��� �9���x����#�v�Lio�������(iF,��Ѝ�v����}T[�$���E��d�>/�o�DZ{Y7Y��X�R�?ۙnQ�Î�f��x5rT��Q��rw%z�6ܫ�p�Đ͋45b������*�G�em���B�;�r�`:��}��!1 ��R.��o+�&���*ؼ9��N�M}�*®��Cs��9��кw�������{m ���~̠���_�c�rwJ�FW���/�PG�ZQ֡�%�I���8�2��d�c�� �fu��e걙���D��aS���D���M��
�E�u2+����-p(�g��:�Y�^�l��gf�쨀���(��n�8�H�G�g*�����x@x 4����wW&A���R'��!��z�h��2���������&�o�#��nػ��KB�V:$]R#��P�	��j�i��V�N�",�+�e��������D��F���4�Bc*¯o��4��Jj��6SZH�R�bی|�����S�W�A<L��d�L]dH}%�I}��(�YDb��f��	���N�0!	tj���s�j�$ohUe��"�ؓ]�;Ԅ��x�x�9�����h ���Oy��W"ֺ���9�ZeL7�ۼ�%-��o# !%Ȝ�3��xUV}�����v�Z�o��x�9`C��;N.���=+J�|9���O�M�N�&-�8�r����<��2Ճs�x��,�!d������O8ɔ9�<<�,��T��:��?)<����E�T��Ɗ�))Hۯ#���}x^a9grz�C;ߥb��1bN��8ɤ}%���T�V�F._�A[~"ѿ?l��'@�o �j�0�o
SkT$s�uͽ]9�f��X!l�P@ ����Q���J86���rE?b��o��� Ŗ�_�w�T_��*�I�Rcz�_���QK�B,�:��x�A�"MqG�X��6Դ�=�(�X lRV��2����dj�y��jf1�خׂE=8b��8D|{o��/6.`
�{֪��f/U��˳tӷS���2Y�r ������pr3��D':���*C����8����)�K�0�P�\��K��Qoy��,Bw�t��b��sNf���j�:��֥��,��$�2n!]`*lTҘ�o���}k��"��D�a������FK�
_Zn7�LQ�*x6tϱ�-,�=����1uP�3{�e:��P��|��^�@���J�5�ls����ώ�,�Zz��bT�1AlfR�x�����E5�ƹ�90Ѯ�EY�-;d�k��B�sPES)-.e�P��a,jolH�3��P�3�~�+u��1�['��oR}�D�N�z<-��#Ւ��h�P�7���"�z���J9m�R}8�Xn�/ h�����wo�ݫ�eZ���W`@��[E6���0B��C׌b��PQfV�Ѡ\�%X���Mq���:�M��,�[~�jOX�w����G������t@��:W��>���Z#�U�é�H���ec��lnp,u�S��M�q�'���a`Ϲ��=��o3ǂ�i;&z�Ý���V������d<a���5�S��"KA4��`M����D<H3e%̷��G-�oؒ]B�&Y?��:(�'�fP�T�G���.�����}1�&���rX�ٖ;� �o �*�� �)Z� �]�nsɧP��젏K=���7��ӿ�
��o���D
z�.{��s��+O^�כ����x���ȿ����ڱ��A�ojQ�WN#��Y�6Ü�+օ�s��
��,����`s.E���^E�"�0�(� ��V� [%x͕�Y{"'��9������<����r ��dt�c���0��g��[v�؀Yj,jZiI�ò2B�I�����9C��n+�S�d%��9YA'c��u8���ﺒL���WU���7����߸D@����0��XHP���:�7P~s=�G�OI10�Rj$�
����T٩p�M�w��ʙ\8�aւ�[�;���Z`KU��E���H�_��P�O(s�#���pD���J�ũ��k41�欸�:��i��Z���� ��,|�j��A��)H��&��"��`E(�]�����;M���B}E8j�cWY��������4�؃o��-`6�5�M���,�^*����㶈,2]����f��:�ٮ����,�^�~��/�H!.`���o��k�U���)���E�,����z�#�{/öW�(i)��BO7g�3����#&��3NKA��Z]U�w]5��\��X���q����*9\�OE�i����Lf�<���-�!�x�V8��L��^p�;��Zg�!���ٚ���\xs����aOǡ%��3��D�D<��mp��F=;WM�6�v.������5<2���s��V��傥�
K��v�D�`r����2g����:Ǘ�c�
�&G8�\D���}U��*#�S����{7�����v��0ѕ��Fa��P�,T�ܫai�{�̨Upu̎�we@b����C%f�7��b�P�����h���G�(�J#`NR���d���[�Ĭ�eJ���'�������o�bݗ�w�.kq�@�1_��S��uM�M��3�
8��O} {5��{�J!���xg�b!��1��NK3�X^ˢ�o�˳sǭ�I)������Ơ�N�����@<��;�Q]�n�_xa����І2���W>��E�M+��r� +��3�v0��S�
r�K�E�pF#Nry�^-���i�q�=%�����!����v�7��Χ�<6�$��2 v�u��@/��SXs\v��8T�W}�m��3�+hܯ�{�?���\�89B6L�A�8W`Ҽ�*�s��MfT�^��FMÆhVý����D�"0&���vf�=�tL���l��v;�ѓ�{`��ǁ��u�~��	�v���e(z������N�!a(�"8X�Öy��el�'�F+^��z�Y��Y/�Wj�M�b�NA�8����|sY�d�Bɱ��e{�`퐵i]챏x���]ͪ^�z��k��������d�{.2kQ�����M�@ӟJ��PkkCcR�5�y��(I� Ν�Y���8.�C1)�}ei}����I��'�nuK�{k��.������/r)����,;*5 ��Y�ݍf��*^k����
/���_
��m\�q0R��aX�ߋ���*�e��g<�B���S.a6�&G�Խ�Ɉ��bV�5�����4/�L�=�B�Q+�.�(�h+S���s�=�SP�:�CȨ�|X�Q�� ��<ml����~_�1�����k��$�1a���rlI�_���+'��l���/����ˣ2�8�˜�Ղ���wpox� d{A���+C7Z��U,AN.��,���\i�]$��M������7�/�f1&��Μ&3�W�|�zCL��w|�{w��3�e=.�VIj��X�hv�p�����3�).����WXs{n�\i:��av�JAM�Dk�j' 葡���`���J��<�<<=m�U�w�N��zL���H{BI�K�}n��˴��L'=o)��/�,����C&_�VŘ~����F	�mS�I<z���+��D����[L�iby|��,�D( �w��������L��h�n�SN����j�.�R�T�[C�b��^��4��mĿ|/8���\��ޘ�x�З�z��:z$1 VJ�����ni&[,@u�>�����/����?J){>�9�e�ҺE���m��a�ki6����D���j.wf����"Ku�����XU؁�t�o�f���kJj�>�Ք���K����g;���3�9��ù�{�@�f�,��b;�ٺL}�/Oda�sG��)����I���i���Qt��Ia�̓#�5ɽ�&�l����$�e}�V��?* �B)��etfGA�^p8�^i1��,���N���7ݦRs1�)3{[��[��F�#�����uAF�@���#8'K��Vae�}K.�0�e7�\��n*�2��8��U���2Ig+=�&�\:��ɉ2���8��]F8��Yc�~�ҥ���φ}v+]��ڨ���5������ ܋���?[���o�����n.�#.o1���%[kj��.L�$}ȼ���-�r,An�@]�mX^�Z��	���-��3u��
)=�cGe��
u�N���f�;�п�4s�vu��z���}ZB�i�b��/�<��p�Iv����qh�P���u���O�D�喝۶���g�G-v���h8���I�n�fE����V�`��JC�h�P��8j�N��^ɼS��f��ř���z�%'�������C��� #d�"5"��+k�+���p��1K��S�$�m��Hiv��q �v�]�������Ķa���-I	N_�fk��h�E&�KL�ǹ$[9�ρ9_�dg���I�~�c��X�����Br�\��ѥ}t�����~u��:�\��3Fd���~�U5�#c]�������rx���s/�p�P;`�35Q����e����{�&���*o;�a
=��OyvL��Q�n���{�^�fWj5�_��Y�u�;b���������ъ��9j�Zg�*5�[vd�K�j���7�֚��`@0�#G�\�^�^�����m����ۓ�2qz�����<1�L�W�D����[h>v�Uj�7��Kv7LA*K!�0;_W��Xt8��=��:gzQt�;<�0Oխ��,���L��	���A�~cӨs�GE�%��3���Fe�l�(��������ǲl��/EV�xh�u�{�zb�yT$+M�����Ѫ�N��Pn�)��$sƓ��O�vd�
N���4��D��j�F �&�(PW�5�/�(h�tb�Ӫ���d��8:ണ�@����i�F5{��L{�@"P��N	�ꀡ��Q���9N��H���m�s��$ D�z�H�n�GP%BX�&�d��1����!q��8��<�����\c��
l{� 0�W�{��;L=0�m�Z� +��	�#�${]d��L��.ʏ7�њ�~/e�O�R�]��̞��5\���wɖ���r�y���.�e�雓�� %dpU��a>3�k"�	`y�e��p��3�Rr��#�-oD�<>0��-���?�.��#y<��X�ݾe��J��`+�⯃y���W���G�L��-!3q%ں����z��bU��X�,��[��Z���:@�JlM/���c�j�8e�WS,���vik?�&V�Ŧcf��x�C-���"�9$q%s�6����z�H��IVK�v�p����E`ڛ3S����'�'@�+sWW���ڳ���)  2އۃ��S�57|x:}/�0㱽�w���9;%P.�W�{�����Yb�>{%�@�Y�z-�r"4���1R�؁2C1Ziy֛W��P��_y�K�5W0�\���5�����E�0R��G�S~���u���{�Ym�D�~��,Mz]Vĥ��U�RZ
�\"�7`.�j1�: �\��3�>���e_RUś`��؏[J#�wS������·�$��PV�)�I�<�@��d ����������%�Ly��>�5'�rc��z5��w�����������a��`Y����+������2摠B�#=�ZңN��G���
n�[�p�pLl�"3���GҪ�\�=�z{�*A2ذ�d�/���p��^�r8��(���``C Zm/�f��߻e�ջ^W!���~���\�����Ϳ�F��۵�y�}~k��7 �<��������n�^^��_�F�g"�"([���o������#:n�<9H�y�m5G��C[�~�\��u���v���i�Xj��'u~�O;���^��>㿇���*��e�$���,�z3�yZ�Z�����TXE	����U�M��'m��Ts�~"�ȕ��ϐu=P��㾓��2��h5n�)���u!%,�9���U%Ĕ"��ZqkX�;��*ؿ�p�)ͣ��N�D:2� l������T]�	����,��~aևP��j��6�Yp�d�ٹ?6�ǵ��\4.8*��M�7�������1�'[v�fEv+�J�]%�,8������7zy�6��#2Z��y<A.�y��������J�ϭ�����A�rW����H�恵r�|/*��u��OJ��ۻ����"�Vf��	��7�k_���i�ʛ� �ڸ1�T��h~��[������!_�<K����$�lڑg���f���.�|�#��R�O��w��v�^և�Y�T��ʍ�je�2��xB��	�-n{�������W�/� +�J�s%��5�}�Ӳ$ul�}8��Į�Q�{y5 ��&��|�l�6h/�"7{�ȈY�*��d.| \�,fHZ���Z�k�e�8�����}�F%Ky{����ݰW;���5˧�Oy��ɳΖU.����~o���*�l��E9�xyKV�ʾ՛������Ym�����p�B}8�I��E��έ2y�]!����@�������	"ĝ�I���Cg��E=[��iqa҂��uvE!����r��Q�4m����i�y�0E���(��^��&h��}C������ۮ8|�B��7y�:6޷������8�o�g^���k����H�7^X=�U������Ce�����u���{��̹e����\�-z����Ko?��{hԋ���7%����BW�-i"�6���u�����{�M�%;��C�8���NgD�N��3���]��vĹ���w1�a<��!!���j؇'�0�:"5�iF�����^C�s��j-q-�Zf�fP#��6�b�<��D6���=ev�I��Z�d�����d7+��C�m~���y<�{�\�}r:D˩,1EQ�2��Ӣ$�)	Y� ��e��)[����M+�-��ӡ�`��6	31�`0��\�"u�ݿ������q�?]�1���~?����,s��BXq��}a�7�W �U۩�rŪ=�V��8޵����8>����wy^�j�w�u�u��Ā��?��Q8�7�7�9�o�3�<ʉ4��!���4��K��>@³l
JkL��nj������K���G��5�J]i,��t�i���b;`�h����Qkq�פp�Z�	oK6�̈P��>+�{�ԩ�?81�XM\�$Oǧ���p�r���� ��$|Md�����_U~F�Gm-N�8t%Z����e㡟�1�x�^��/����nY��:����/~G"b�L<)��O�e�]�<= �2�)#m�F����X��]������oN��g��\oG���w��6����-���6̾ن!��G����V����&���Y��QF��w��	[��a�ؠ�W@��7��E��܁=o�*\9�$��F�_�8~s��%)��/-1�M���sY��=�����~�1� _����K���w�]��Nߥ�вu@ٜ#���]�	軔����\�F�P��B�s3q���|-����о_���� ��^�Cl�lї˅���|��^�\�u�Xq�=Q�M�D}�K�W ��V���K_A߅�%�lUЗ8ޞoկ�c����
U���k�+�o�Wʨ�;��)-,����Wo#կ�F�u��w���~�']�.O�:��b/؃�G5?������b4ӛ�eH���qGoWN��D)׬�ެl�V9[ן�e�Gy��/��hL�)�O��X�>ew]��������k��dII+}�A�ZpMJ������<1��>�q2��-�k<�	-|�w~0>>y��ҡk��5z�M���E�1vQ�f&�u�1�veD�> q?M���27��0���2_�z��UȡI�#��]���m*]v.h��@cl��WZ�4$�� �挴*���XVը~��w/y�{�?��>5�^�{Gb�Tm�����@/ѡ���h�����=��;<_�!Pnr�.����L����C���Fn����-�Ĵ�cy���w�:{еIs�E����![2B�$jNP�t���7h�O�?��"Ϧj|�}���z+���z�Nv���Aw2�G�r䘩8
�t2�rGSu�%��z�^�q���H�fq($%gt싍�]�o����Iy0/ډ'8�M�\�3�.�N�z}��јc��{�IiY����m���UZ;�d�Z�k��H�}�I�9���r����3��NF�2�C������]�a5U�!���� �n�Ӻ/��ເ�z�)ǻ%b��V�E��!��Ul����Wz�4���9��mNۀ����づ/�+�}s�4;�n$�Χ-��ؑ�J���ʡr,��o��ZN��=��n��s��_O�]�L;���Y��g�΅�$�,��M��zx�n��MjD���XSVRI�m�x�*Q��t�,����s�=;�c��sKzx���c�Oy���9ͱw+k�ʷ�Iq����o�>��G$8�vw[�S�dj���i�����\G߅׸F��c-V��a���ĔD��,��ͱ��w�Nj{�:�y�z*��j����y��o�N�ℭ@�c+�{��$���8S<bSMO�|Hݙi��}WAʢ�oB���:���]4�����D����~X��7��.��;)���;34�T{7���ɇ�?�����W���(�)�N5=#�2��1ʟ1����w��5�I�9�n[Ny|�]��X� !t6�!��JbYM�*B��%��n�}���ܽ/�d�I�S�m��U�8~�H��S�P��F��e�X0�잓����OZF��dOPl$�xݣ1^��+?�z1Wu����6H�Ϊe�ױ�.,*Z��K�v�|4���L�$I%Y�imj�\�!�>��[9��1�|�dIѡf�dʃ���a0)m���08�V�>�33��S3�ĕE<�5U��&,"�;�vX{DP�������InR�g��K�ٿW1���/�(��FF�d�ʚE��CO�e�_3#p*��tt2s����.!R+l��b�UP�_D}^��T�	�i�fk��Tg�Y~�|W)=\� >�%�o��~n��<��I��������B���%O���+��d�N2-��{Y�d
B��M�e���]���h�EUX8�2�$��7�W��+���w0�1je�W�{�#ۃ��[4�Fy��*�`ř��H%]�u��A�����^Ad�6N���^
Ew'U��f�:��$�h�E�z�!�Yb�ES�j�`N
��B<x�{8v�rC��j[���33=]ባ\��)�QC��v�/HR�T��Jm�ma�W��`�=����Blx�]�g�J�Cb���V`��-�D��xo�J�	93�[(��R%0�Wx��
5��2�E�'Do1�K���?��5 �ٙpy�u2��y��$3����v�A��7���B���V'� �> n�=�Zjb<�?ڗ{�/�>_cWAq�M?���:S׶9��t������"�S�D�N_��~R�,X�|fft�,	�/�݁�2)�|daoI�ߑ�1�� 5kx}�A��!�l�K�#�� �U��N�A������$�#s����?�z���m�yn�� �\���	���Ī��r:X+�/��"�j&F����y�ow�U�g�G?
G�Oa��8PKt���	ƙ�����^=�u���|�v%��n��mP��}���h�c�����.��v[;��#��>�=��*Q(g5�3j,J����ىK������n���s�2_~�a8a5�ϡ�o����Puy�̫���d�ۏ��T�-ܹ��G-�ǵ:��"K��]o�&�/8E��T��O�WW
��"�C��_���x�Z�%�,!�!޲�Qn�i���=��>fR>C�,�� ��P���(��ns��u��2�q�� <Yo��PTtl�`��q�E���	lgݲٔ��  {B��R.q�GF�E�������qLZ�J�ڡ�3�k��۱q��0�f�E�@�#����BH#NG"���E��:���")��	�ai"�N�.��T���� � ��G ��VY�7�Ќ�V"M�	1�ޟ�_�|�U�{v��P,=-ݖ�+[�0~���I��0v�N�+�_�>�I��+����Bܞ�ۤ���K�Լ�m���~���D��z�3d��&$��HplI�Y}3Ϯ�N�6�`^hH�,h��)s5�7�x�Ğ�=�f������^C"�o=�l�;��Q��:��s�" ��o.ȨQ�.�%���یh1R�n�Ffxn~,j����Mdz
����J��4e
P۠�,��7yi�^�ɑv{��iy&��n�"��{?9�&������㋗��:��c�.���ne-x�D�"�B�Ǻ�s�UB�P�r��A%�ᡃF�6��d��	����;�^�S{�����M��r^���53i���L�s�RH[����O�ׄ�O�q����2hĽ��MVE�ȣ҆v��+�/����~�k1���"8)�H����1K$~~���?���!�Zm�u`��_w���"�,�M87�5���a E�
�7��6Jp�`�g���|?Q:^��aE����r���C��i���0�*�3Ŭ�e��z0fv�a *��\-m76ڧM�:�)?���\쏁�4�Zv_��Gw��9w�ֆ@������w\ߴ7�ĝ`qձ�U���� �i��?��7��� ��%=�>�q�Ք��t��X�rX��&|��g������>/^�jcʮ{*9���Gv&�O��R}@Z�{�]�m�E�Z�=�X�y}jql�J��R�@���!�f	e��U�O}�����:�%��O�h� d��r3NŶL���̟Q� r4�^�:�uO��9hu,E�hK
���!����s�%`I���� �]I��f.�|���d\p����:[�o�s��Zo/��=.��Xձ� ��t��7�%{��N�S�)��]����$z�٥$cH�@Ћ�P��`���A��Sg�]��.�Ҙ�R2�RD��3S��Yn}ei��肟�C�9K�Jٳ��̫c%��a�{��n��ؐ�ϟ��c� ��7�oH�>��{�vq�-�_�����B�sQԎ
Y����n۹�!��k<�]2k�|ui����kqRچ��)�k�o�Eb8���4]��Ǭ	R�/�
4r�5�ه8��LT�AB����A��2�A��&�����(��G�)s������_�f�����L���͸��=P���ex�o���@hh�qv︺���mV�se딹@��t��b�v�x�u��1����I ����\�U �T!2vJ	� �b��$*�OޝPIC)��#�Y�FT2�$٣1����He��v��}���1~|�����n�#�D�Ő��E���#�۰
�u����C�v���j�.�{����g�@)��!*�[�|�kK���i�ӌO��'x(�L��N� 0����vnʒ��|��X���,�Wɜ��Z�L�Sk�	���s\���}�(��*R���iC	���s�oT�궪-s#YN�K�h�ެ���na��p�{�,��v%̾2����!�ç���ચ5�K�!j��C��-�Ý֮����C��l�VN�zTO��PE�^��Hʲ��U�a�+��v
(iB%"��?�FC�!�;�-��k��a�;�FSuf�#7��EG/_���A����Q'x���s`NU�L1��`�LZ�y�^V�w_���t���o�fT�
�m�Hgi��z �K�tJN��Fyfp�7
��%��v����`������Xu��]�܋�rz�(b�[�}JY�AZ��^� �z�����,�o�di�����ODl,�?f:�CTO��!0�� >f�u�/�A�̈�Ӡ�a?6���Ҿ����hE��	)�fͿ��[z2q�-��Ƥb1L-�hN��[�xh�E��J;� �y�mF�QU���..�/C��,�{�w����-o�|�"�8�
�hۚ��  ����AϵM�}�|��z.�t�2�sd.�!L����Y^X�$�Fo&*6l��]o����7������x�Oߕ��o�.���)"�'VR}/h8��)���Z������I��<�[��e��T`���c����?˞Q��7�i�o�M��p!8VM��/0�~j����R��QA�* h@GH�9�g���ʢ�W���^*��A���#�ۛ٠�[B��z����Yڇ�(��o�g �3�6.q}�is{�����TH{�v�A��B.e_�X[��F�u�v$WQ�-I��M��c���e���ԧ$�4�����l�RF	�:��?6��Z]kF}�<�lW��̵��NX�U���ow�B4��g�23gj%C���6��]�!��'�x�l�$�l�ոv�▶���W�~;�k�`gf��٩��A�A�������R�É�)3���R[Qs����}CȨ�b��v�3�Π����:3V�j��]�Av4*�f��1�\0�_`쒓7�~������$'!j�)���z�>�&O�đ���b�Z¹/t�Rs��>9��]�<���e]���o��
�h��<a����U1}��I�m��x��������ǃ�2����o��d���m��E��ֻ���s0
_C�J*�����^+Ց�uy����ټ�cW�e�M�kj�Kk���Hk�2�L�+��w���B6�z��(��>G~)`�~��t�z���UO�.�aH��_��P&_zO��:�|����:�$��6ysH �[R�Rv`D��W��G��_�����>1��Nk��?�Mi��DT�m�C���-y���3k���6l]"=���!qV[�KR/-��)��Y�)WZ7�ϩk�"�x�A��ȡ?�p3��̠E'F5PX���mz�~�4��O��AD{���_� �mʐ����:���a��E^����L��i�}�����v�9OI-nH�׋�k��W+�܁��f�=%���e��=%�qB����V���DK�F�@������)��ݬ���M�5܀��M��v�̃v�v����L��=�n`8��t���0�-:������h���ȵc}9�bM��L�+��O�TjUpő��,�}�$�/AU���4��B6����>H�c��\���W4�W�>��z�~�^�q8��n�?-�3eqs�߉S�#�!O|7<��>�T%h4ι���zCY�#��k��O;F��>>�-I����?�e�|�^� �;��������/�{['zD9,<�s
�}�Tr�ʡ4�Xo����b�$� �Cn+��'C5�������ќz���4v�F�k��J����Ʀ��0��z�t҄k��d����-P�~�G�c���,̇�¹��)�HA� ���a�7��m^j�
6�Lǳ,*���=r�b�C��	HVc\M!Gbf7¢" ��{����[Y�� }ZB����D=�훠)����(�d���x#3�5A�*�ˀ�N�Y�jrўO��q����%[bȁQV�o2��RU�ӂbTĭZ��:կRꛘ�Z=ɛ�ό)�Uu۷p?��Tig[ �aiW7o����n�d�P�p�If�Y�6x�}�
��3��A��}2�^-�?]2�6Li���}����SL:��-c^׾�9~S��gNr�&���I}�l��ô�)��(���踵�6Z�4�H��.j�nMt՝f9��J���$w2�h������<�������;$���fٴӓ"����f=?�hG�9j�.�%sWvׂYz>���	��l[�U����0��X9���~�EC$��� j�Hku���}}1��S��۬Z��d%�E^]���Jgңz���j�f�1,�=�b���dĔuoj�MN9��L�I|���	��WC�G�ҖeL�R�t;:P�ϱ�;�PX�d�j�����3�ֲ�{5�h�7GQ��,sm�g���ݷ�mB�}�4�l �Ͷ�<�Pu�� �]M��x���|i�D-����.�C��bs�����+SB�}!G(�W�$<�������h���`�3��U��~�u�a�����6��e{t�"��ꨊ�M<|��{~�??�'=|\��VY��P�(z� a��q<0^(�"�~sA�I��p��L}����?����,�H2v�2H��]��z�u�����L��OAf��H{w�,{\��E�����E�B���ق�\�	�q3�a6-�M�o=<��!����p�	���^�<�z��@����1��hdy'�1+�ar�X�	u�zO���̬���j��!���a���s��:�V��i{һ�PR�R;MD��	��M��L��:K�M�[�&(���8�f��}����,���a;��x_;��_�&&C+�'H{�4�j�N��,FZ2Yyjf���/��p�dI�u�����^��]H*`�x��:�Ȗ��_b�e{^+>����F��O�n���ݤ�������"H7������c��s�Mhi��e}��b���RCD<�0kyo��a��PD�����s���g�}� ������ْ�b��~ ��|�I��p�8�KZ_��ۡt C�i_'�G�P!�A����>p[,24�z*u�$��ޓ�꫟��ڹ�c�]HY��%_�T�6�e���/da����qܑ�V�e�i�;�:Y<�5���΂� ���-`�=�������M�gi�����qx�5���W��Y�ϔz�;?<����㲎8]�!$�_��af+8a�T�%��1�A����=���
b4����~�<�q��Enz@���H�&^I�s!�z�^)��ؠ���,.4p���f�[G��X`q��~�@|۩q��jkykv"O�\)��{�u�Ȯ��|r��rz��@z��i�G�&��-���;)<��p�{���UZ��IFQa����\��忌1�a�y)��7� �=���\�˶�d��Ƨ���]- �?x�}ȹӻ\oHX\���+��\Wt���%?�1����2�%a����͖l5y���b��ׅ6�X6k�%5���ʺh�nY��Y���8/�lr9¨я�8���o�3�P�� �sY���fI��8	�	+N�}��
���?�v���`o��Dk)� ,�ik6��?˸����
�ٕ03��lo�)/��B��ĭL�hO�|���)��Qk4?�Z��=I��Z�����Vʒ�� w��j���~zCƉ��R��lX���%J���ؒ�5>�ަ���|�I��z�؛�2P������sa�C������o=.��mы�� �O���&�鄾��=<���o���� (w�.V'��\:9յ�2"�l�	&�\�.8�7��1��%���$������q��΄��}?�	�ϿmmU8\s�xgVٟ�5���':-�Z=���})OA؁��DvK�6�=w�����J=H�PL�T�3���Щ�SOw�,!�9�%Im����]��[�q՞7�2�Q�0�k�xS�t��)z�)�v�bKHR�"0���7��[9E��#�v,թ�?r�P;h��bz��F�hߜmS�4��¦��ܺoRWp�_���г.G {mP���u��6��J�-����z����1���%fF��+wZ���c�]}�v�Tz�M���R�����b:�*B�m]�s��D:~5���kw	�mփ�ɑ���"�5' �8�*�#� ���ayB��>�&�>�47Y��y�n|��9�,
��*���!)z��2�4FrjX6_M0���C�#�`��d�Ӎ��<��e0��#?�:��.�?,(�X��N^�t�QhYM\*���p�x$Yl�c>�u�4ְ�z
(T쿨5�c	=��W�2̔��x;�����!{SYo�Gfщ�[��P6���|�rU�i�N��z�6�����h��I�]�%&m��������y�P��Y����0�Z Kc����|x�_"�VU��R��f�|��������}\Q�O�\�qY���L�1�v�
m>�)	��h�2�JٰJ��Lu����!�M][L��.��t�LhU8��=İz��ͫ �e;I �l�ԶX°F f�����l��Az�6��8u���A�0ZF��u�Ww,�����Q�$l��~5�_��rPQ;�Xq�x�,�1��%��~F�C�0���!,�Z������ʑL֮��n�P�m�m�̩�k� dPܗ]�ko��Ӂ� �Q Z�j'���UDs��ŧ@�>.��Iv �+��lMy:�����4
�Φ���D���}�ч��+�5�*B^�+^5�HDy�rF�陋�/���Vh�.>=F�W��Z�ُ9�g��]w0WM;�i�M���_`��F�S/@<&/���$�`��vk�.�{�Xh�߾%�L����\�Th�آ��xu(jK�Ȳ����r������R�����I����Ч]�����h5������~�� 	ht��װ[��$r@�XES���b�y#�QmП;Me���#t���Y�g�b��8!	�[��M-S5֮�n.I�P^W;�<46������Z�gJ��G��̓U�dwS��RROW�컺R`
+N+�i�%A57�t�k��"��ϸ� �������xu�^���eC��n, �1I����י�Hrq��2/J�A�W�����@�y�WѩQ�{}(�o;/���;Bˑ�٬ѳ�?,�u��g!8~}�7I� x��s@w��W�%�����܊��.dU�Y@��T�ߦ/��ި�)�v(�jl%�+�
A+-��~Z� no��Q�vq�i�v(4}�d�㫯�ұ��xX�b/�FA��}wP2$~�"ĕ���x5�^��yg ����dNڀ#�jUG��pcB����K`����6(!��C e��:�<n��\�6t�M��V:>��)���Y��k�榺;d
�~z��'-����;���Z��O��A��S�T�D�&��F�X�Ҳ���֧-��
���d�����**�|u/��o	����zT��7�RQ���j�ײz}�o�y�>Х�˶��� r�&!�ɬ]Y��	�6[w�� ��?iN��ڊ���z��ͺD�� ���#G}�͗�UG����y�[��E�y�/���sߪH����2��1�l���V���Ȟ?M�<��VhNC�̝1�;������PC�US%��S�i�j��w3����� ��( ���[��J\���OFO0�3��c���`��Y/�������AC��B����S0��]�(��7KNULڿ�>�U�l?-�{nZ�g%zv;XM�����]�����(����*���o�@ƀ����?��d9/��o]�~W��LEk]��(�%�Λj�'5ib�IiO����Pg�f�h˧ddY븝ˉ�i[�Q������q����G���Fz��16���߁��
�K��Ȯk�w�9U/~w@�XXJI�Oux8��g���� �eVg��4�$pvHA�?/�����i�����4���0W@���Zj{}Vj�V����sq������уW|)�`O �l�.to����dZ^�����[W�N�pe����?{R�n�>%N�$3"�J���Ҵ�)��c��A�#&%ZbjGU�H/k���U�x�Lg9L)=|��O�E(�i����V��t��%$oV&q���P���3�0��в�m��%bY�}e,8���.��S~.�%Y,T������Ao�K�&L�C�9L�ݣd���S�|TK�%�޸�9<���7M�8f�è4Ԁ�}�;���oyX���zCL �3�~�j�]#C�;Sm�H���:|DuCI@*�^�7�m78�m�����r.���+VH��� t��-�˦����>�,��gi����g��A	E}�qj���ҩpcl"�N#�Ks���s(0���P�dm��w3����f�`�t������/,5�f��o�2;��ʘ}��FI,�(oV�d$̈MeW�*�<C�Wˠ'%*P���_����u��Zb���g�
�L�t���?�P� ���WL����m���{c�]%��-n���5]�/�(nOѨf����d�oO�?#���,Ma�cque}E���a`��픣4W�ϲػ�C;y+�]z��<���z���94�p x�b �Mc9��~>uH�-D/����|hyv�l��f /� �5�^<Λّǿ�����F����x8�Z*|�E�!���"j2;���s����������~�ku������lHN.��0�{���4����)Y��C�!����9Ⱥ �`#t�/B�"��U3O,��]�ɰ�x!� vGkʕ���އ�שHǔo@Ke�ga���a'~*��Ě������7�#؇��'u/��W�:2�=������ă_<u(��c�>��'ypf�"$o������i���`!�_�{8ۚ�ԗ�v��dE�
�Y�@m+u�m����ͼi�����nm":d�Uz?s�e���Թt0�ҘD)�F�u3�#�4���[���\,�c�u�X�H��P*��`�����WƄ�w�6��n��,�7aY����tf�)}@xt���e
~_<�n�>u����{�~��BnyY=F[�f�[�=1OQёl49Qr�q����G�0J��Q�}�~z��`_{!/�ă*����47 u@�g��֠��؈�D�S��BcV���@W���剟 �}=��U�{�*�,A�V;�ց������+���O�]t�F�pFL�d:� �5uc w��&$�< ]Y/A�H@t�[
\}��B������h�~�=�1H=��Q/���V6���9�6Զ#�D5���z�ű�:VZw�R�Z������s1��.z"7UWa��F��)Cn���E���ϔ�Hp�j ���q:b���E~�?an��������8�LGB/M񧏺��ܦ��M�����ol�O.��cRR#����گ���)̤�,�tS1���W�u6��� ��]��&R�z���_�~�����)���)w�.����̴c�*j4V�g
�� �����f��Om�6g��E�,;�O�Z���� X��[^��7R���. �*�t_�c�#9Z���ԧ0p���+6���)��N�H�s ���c!A�O���~jM�BDά��r�	x���Qv�U�뭰�U���ڨ�A2�㫮lo�P�s7�g�Th����Xj|���Mh# -�"�?'��󍪾v�v�}k
~��~�懶�^F|���xYz2XC�!��o��u4�� ��o��u��u��|p���\�f���Z�~z|$����{�?�?p��"6k>X�����?>�ӺK���a����p?�~h�?\+>"�P�R�K�.U�y}���_����V�D����������,��h?J~E~(��s��շ��\+*��z��֏�$�L6>P1U�}��K}Z����w�
^�lJ_�����S�K2� ��e����Ty���|킩�L�9f��q�a�vi#z��*4�Q�����i���e���5��C?�-`�$��gL����A���w���q��p��Nl�P8#���;n����B	~wX�Pfm)�G<���6�Lx�E0���D�-��)��j�b/���UZY͞:/�������6^�XFCAz��&�Om��ε����D�aY�2����K΂�c^��=�I��{���K>�v��-.l\V@�bS��-��@���I���/m�?�.w
	 ��)�J�������$���8�/'�hsʪ���Vk�ƮCW]5��� ���ھx����X�-궉���}�K
�g�RSkܯ�M�$�5�r��Aa��1Z��/�
,�w� ���K��5�����_5�����9o&��LK=�g_�i��X�ᒶ��ӇQ�D�Mx��ޜ��-�^Ѯ�{�[��:�+c�U|�l�?]��?Up9Gm�����y�i�)�0N*���e6�cX�}G��7dF0�%�g-��ñ�vh	���>�\�׿������lv𻜖�!v~�*�S���\8$�T�0�����ս�Sm[E#sE:��N��&���u���m��{*I^o�ק��V�]|�tĞ�����5�7.�
��
DP�sG��R(&�<L�}p��&:�4���Dܮees��ݳ�"!���D�-������DR�{{��} �E'��R`�r^YT���V�l�Y`4�܅��a
?D�ȡ����l}O��)�����U�`�Mw����^_��B#l+4��u#Df�F����(��6�	v������\ԇ���p ����i�m7��sxXqʹ��{Dw����j�/�^�<L��j)e���Z��^i[�w ��uF����X��|��kZ>�.� ��i�Zx�߶A�} �� ��D���[I���xZ��u�V,V���@JI�^����=�y���O��� ;j�J��YS.:�->���@U,V�w���5g_C��Co��Q��4�װ��$߬Į�ٌ�G����b�،���6L7I;pD�Ξ�Se���/�z�`�l�l)�&қCmO2Ej ����l ���rњ����2߫q��/A��f�b�U^�a�>���|���z>�7�qr�TLm7�N]҄�@/�y�2\E?�'���I��v׷A+�$�M`�������*��]����@}l���/����l�j*��8N���b��^���0�p)k�sY
��ο�{����Y��zq���_�|q�h�Z��ϰ	}��l�?߳'��;��_�_�-�u�]ge�|����8[s�/� �3<b��s���PK   O��X����(w  +�  /   images/42266fcd-641e-4cfa-a619-b442e1b7bf10.png�|wPSo�.,�X�( �KT����t�C(�;(�Ho��;�)���Mi���йI�}�9ws�Ν��a�	�d�k�{�g=�Zk�PMu�kT�Tה^>ע��(HAqf����贂��/�߽�s��0T �;s��39
��)��r@ϴթ��@�c��~^�Sy�m�?H�����@����&%`������;��Ɩ����*.#9οdC6��񕭖Ĉ�P��?Y³�T��^Ե�y���ݑb�ћ���������.{�?ާ��<��7o$�'������������g���+S�*�%+���9v�G���4t,�
�I�@A8=(��#�2ڑ���,�����u-��k�E�Cps%�%]-
ϐ��G]����[�?ffL��#"�yd����gP�==���U�c��\�}�?u�IN�OIIy����2�\̗�GOWW�����k;�-�YϤm4b����}��Y*��h�+�e��/�tP�i.Ӕ�����#�϶H�N"�ii�H=�).�%Z����\��� ӿ�F���N���/� t����Z��N_�~���ӝ�hY�4<<:w��Gxx8D�J����ML����#O��	A��ҥXm��k+���|�*�[c1s�Qf�C	���e����~s��oZ�/	�ǥ��{����������rw�b�0�C�t#>#�����p�1��|1�8��;����Y��h]�/��2����$�i̍=��3$�{����7�����ܩݖ�%��}W<2��ɔ��І������q-ԕ�k����[-����5(���Μ���h)� �7H榤 ._�m*�T9!)���l5Fl��gR���

�_#�tw�}�Y��>=:�9��)�_O����`m�q�vM��R��S�t�8���������*g2N=�-ʔ˲↩�ު7��ˊk�g���\�j��W�7,%����L��ض��h��	�m��V���O�����_�،����^�,�7�uKK���Ʌo�pq���Ù�� �5=4�����jɩDs�!�Yݜ�Y���b���nx�����s�g[o�3�6
����?��g���;wq[�X�|�.a�Kn����{�>p����z����� ԧk�Jo4c���;���P&÷W��\`⾻a�[�)��b����FFӃN����?���Ó@TA�����]��!��%����v��^�����K�j<��/e���nSI��{��T�o��x�{�:u��7��_vb��,":��5���,v��VKN�ê������xZ~��s^{�z9U5)de/�	bQ���UmB�Tc��H����Y���{�Ԯ����,7����;�c�����:a�i�R��I�2�^�2Jq���)++K�P�ـA�MIv9U�@����E��#�6]��8��GHڝ�X��t�1�A�ڏhy۱�7�!��8�|�jiG��:_)�t��o55i5��� �*����G����cXO��[�W�_���+?nph���k핻:i��p���5dɆz��W�@qX�����|�c묋]��S3���Ɇ�4�W�<�����kj�nrg�}�h����_t�N�D�=�[15�Ҭi���cm�^��v5*ύXe����U�u���)���)�lPCP������Cz�w;W��d�/:��+۾O{�����5Y@r�,l��פ��7jK(^0��'�^wm�k��r�������_^F�z�R����1�`@�{��^��ט�����ǻ� V4}��K�6�����cSͬp@:E׆Q�Z9N80~�P�NO�����V�� ��;~���#<	��e@ɮ� =���zo�W��L�SE�2"j_;��g,�m�+��i��grg>2�ޣ�dF��1��O]�l���&^�H ڨ�S/E=|He�/"�}�X�"kTލ#�R����l�:,c�
/��"M����٤Y:s�I6?����!P�#�9���ˢ�tE�Z���cu�ZV�L����'u�f�R��״�el�y�}x��?������"����c�MjMgϳ]sHL��=ҪaNO�
7& ??n��`@��F��F���r����W�{6�G"�8�snSѾH�f��1��4�a��#�'�0�u����/�.::�Z��R��6�
g��=!s|5���t{��2��R>���M�VZ����>�� �M<���=d!�b���ʐ}�����Q�4�_W~(-m�	�C/=�}U,����u�����=����Ҩ8'
oz83�y�z����H@�ˢ/��;�ALɩ|}��n��y�wꍑ�xj8�[���u�H�{��;��7���ԡq(��]v���X��ʺ�c��٦�B�^.ݸ��o��dO,��Ua٩�2���}br�3B ���&D�h���������G&�=^Z�@�C�[�o>&u�g�:V�9�m|���Ewt��Q��҅�b@�m-�6��l����}���&$�p��=�zq�<�:w��+ ��������[��'٥�+BZ%����h����i?
�>��ɷʮN
S�`Я� 1ܿ�� ����cޢ克�=AS�d�"qz��3�h���͹����̷M�,���_�<^%L{��"��l�A�/,v�,��_���M�8�"�f�2m�V6:���*�����3�))Qz�{�`��%�!�A�;D���G��c�w.�{�9���csz�7�.W��Y���;��B��`��zMp*�H�;F������t�?�s,�C���-e�z�A++-P�3����7XĪ���~�l�F��g\}���"���î��Q�l�Ԙ�T�kǇW�h^�����y%��13>bZ������C@oݼ5�$�cr��ks3{�Փ(��Z��dֹ�]Ѽ7�������Qe@���:�� ��/n+���	�����jXD]vxU�^�&�00>�ѹj?��۱�n����"7�l^ٙ�-�� "����+G�ϩ$|q������%-�e�� r��6#�U\�����m�F)G�e�*۵��*�u�Tc��#Ϻk�Ӵ��&^�E�g/��I��-F)1�z�����ί���c�|���vl@�]񍹢���1��a�e\����i�F`՛%�R.Փ��DȞUo���R�k�e����v��I�e�7��:��C�=D���{�f|yV��TM��.��E+���<m�P�)I\G���aoh�K�������L�U�n��/��Z�|U�&�[C��&�C�8��yǠ�t��H�
I���WSfn<�)�^�v�?�e�6�ļ��ã#���-|��D�1�I�3E�y�����D�NI+O.e;6U浺n�/ ck��S�XEt� �Ҽ��Xla�cf#@̾%N"Qע�MR7��^~�Qa����1���c�ny��TM��`lTZO����z��f���G�jȈm�,j��Y�)<e!ȵ��:���jDt{�e95K(���Q��z|��N�\T #�#�פ�q��s�޿ٸ�����Q(��߭�ފ�k_���=}�k�l���JҎ��M�U�D@��r��c��nk����2&���o˽o��K���<��4�ٳ��� /Х���߷e@�0�"�2���4�<@�G�� ��ؓ�0���Uȣ���v�EǨ.a��~�-]-D��`�fAL8�������aUr^s�B���R�a1?vv��3;6���x"�P�]�o{��풴�%78v�En�(]�8�y|�l�FP	�nfE�ǡ&ʵ}2N.�C���M�&���N$
z��
wq^0u=$�-�*l6	�n�lj<�o\��]�������c��&<j0��c,A�a��p�cٓR���#@M������up�7�f��@U��,J�|��I&L�W�S#3��ha�~��p�|��H1�2��݊��OivV4�`�D)g��8#��w�����}  �V� ���T�ݑr��F0}�������p�eW���=�: *�QK^�.ϖ��l6�G���(f�g
i���#�U���uNq��
ڱ{�Ƚ�ЃW^PG�D"T+�s���������2pD3��@��c͋l�]���b��T*�����߻��.�2#���"MRO^�4�o��hQҘ��";�x��͛j<C�,-m��0����m�+��9{���-֍����4%�Ia���J���Ƭ��,[���_f�lG��D�n%pYC|���>3Yg<9�Ey->CgO����|$�7����R��B:����ˋ���l���D��aV֗�Lf���?�����hd��@G��}o���������|k.��Z�����Dd�a����1< ���#���[:^�]5��h
ɨ�"V�����#��h�ɶ�AFTl_��«HQl�}�i;��o�m��j��b�N�z���Ѧ���t�2]�ĥ��r#x�J�H��*�V�.�EŉJo��߯,�����
�O���~�:h�ie���+�Q�1�Q�O��W��x��>Q��Y�����+�t����h�n��כB���k���M��(`1�n��P|�z�P��4=��H�}����)�	N����0#�8ݫބeob;YSܪ�q�JZ�}�o�⫔2�z���-����K�
wﰆ��	(�Vy)1�b����j?��E�h�V�q�����b�^,6�[XtVĈn���]��/O�#W~��:&�'��Q��J�(��qI����������1�µ|�e,��B�,g��lQ����6X�~�r�:!o۵��]��Q�o���@s@~��jC��V�l���̛�g6���v��LO�n�9F�y����c-���k �R��ŀ���b���ٴ��'��˶��3������������6f�2氿h�7Q5�ÊMbY���]�3�����Z��Q&�O��K�-��<�=!�BӁ m}ؚ]�l�r�\Ṛc:���
�D}N���U�>�<Z=���Ũ\��o�0�t 
@n�o���l����X����w�,����
�CӿPqs����$�Y�"�r��m4�G�r�����~=��ب~8�n��DU�x���/2j�<6�Y�	�GG��H�f�|�\��̇��ՠ���0Ҽ�.6�m!�����l�^m�$��}�Ww�9h���a��J��@�$���뼴��l�C�J����d/��e�>3?^) x���M��%52k.��t�\����t���kS���W ��F��2���DpR��T��'�d�p�f���� �e���a�g�O�յ�*�y���*i�w �^�(!k���x�TQ˚��$�}�8�]�L���L�+�GN!�RR`�����pۯ�5��qOn�Ϟ!F���b��>7��i���xShl0~В��D�Ȫ"���iR���;���15"�þ�(�u��*F+7�#H��:��CI����eF>ܺ�Q��e2T:XJ㿪Ljy.D�h��ujyW���kϛz��DX��Wo@�Lϝ)\x�{z,�U�B�VV�Ȗ!��`)�0C����9��ii( ++������uƙ��t�Qȃ�_��I;�Qna��\H��/���A�O{�9aX��9��(>�F>~|9U��`���Pv��7fs�'�2�7���.2TW�s>��D���d&�	�U�+d�o�{�(F�p��&9�1z��G#�cuĽ�%Es�OJ�E	o *٠F�۽�5a����r°M�h�}6A�P	`ץO�,�������(��m�Bxc]'m���W ���!���݃=�wD���U���Rm.�U"�5�_����WꇷP�g���[�<�Y��	�jg��i��Jtn�t�,��#%TO�h�
��h�˗��H-����`�_�L>�a6��rR!ő�6��|�����d������
R�tC骗#/H,떾Y	��Yב�Y��k_B��U����ի�)>>]�
T�X�@n�G
V<�t�!1��E��1:�?
��H�W��/W�z��%�/��&.&eyW�%(�!��)с#������f�
J�-) �8���Q�S�E.*2{`ݘz�"Ea�{x�bQy�h��J�os�q�(U�4��|�X���1��&c�U|���V��f�p����kJ'�ۻ��������>��܌�n{M4�B-|,��������Ђ���*�_}R�N��wG��C�b�E��A�?��m.�(�:/�X#
�c��I��B'���+����cb���&1�%=���n����kt����.Uf�uT&ڑ�c9�i�Y�]�7����������p�;,�C��:���* ��m�a4���� h?�s�.9 [�j	ix�v�k�Te�y൷���mU��S�L�8^�,�VS��Y��ky!sا~��}ڨCߢ��5@����#����f��hj�1��������O1l���蠓��L z��ge�����Ή�Is���~�bp߱��|A�Ll�՜nk�י[���:��z�㥶#����B���'�ʨ.m�`!%�M\����a��W�<��:��rH({A����Bv�1(k��vo�GI�I�,��U/�U ���#���ILl����&YE+{�|
'�ᰱ����2�Z�?�I���/�j	o"�f�[;n�|���Oײ:���4���kX�Tt'��B�BǵTs�` י�I��r�u�W��X֦�J�ݖ�T��$=�T�,{���a�WT���5�'O��J�������\M_iY�9�}|���G�9=��M�\���hw�p��������զ�	B��4_�5��� ���N#r��'UoS�RP�b����!��cs/���m���T���G���zz����[�}�&g�v��c�P��Gc�e�C�y� 7e�t�<���!� ?~��5�q�>�zF���{P������h5ns�0��h�I@��ߝ��p�g  e�7��~[�U�,������F��#���j��0����ְp�2ouD:1p�o+�i�3zܰ�Bc�G�h��e+*�f$!_��Gv@��ъ����"�Y�:�O��﨨��|����3#�c���Q��{�Zll,�fny�	|Ks�	����+��&1�e�j���J=V����;�,F_�FLnBQ�"�{o_wԻ�y!���-)S��s1�|��39IMy`�n��G�$]IyT_w��Y���Ⱥ��H�hi%�7\�5�������i�u1��-+�,��Mx�1��`y<��*q�M����3#w���6�Bk�zm��A3��V�ۚ��-��Nn��W��|/�)9�Z�����C-�] :E�b0���S�Htq�G�ʽ�Ws��yTB=��J�Z�� �<D|�o�Wqp�Q�wo�Ņw�Fvk��BO$� �珎y��ER>��z��^n��=`6�W�\gU�ufZV��˅��g}�ɖ����W�����c�����isv����fdqQ� U�J��V�����t����ƫ
4Gp��Hy7�G��!��zX���0�Y�e��ڬ�	�̭&]�h�^wo��ʳAAy>�Y\�D��ڧ��=�?�6d�5�?s�E��&c!��F�u����ʝfա����{S�W�i�c�K��]�������j���kG�5�B�S�\}B�~���(�Ư:�[����%%��������6�5W��.]���5���먥��׮�W�����]�P�R�j��t�]��V�|Y8Zjx�~�F�x��A�?��F.�}s�o�5���<��⡫��K{���Q����f2�dO��f�O��)�M���X�Vs$7��|���QN% �)��d�@;����i�1c��2tD�6G��ԏ��s�z�j�ݺ�Ҿ\�y���(��Ħ�"�:Q�Q���3�^1��gy�^�vu8����E���?�%�Q ��D�29(�*��o���f��yJɣ�B���o�~���RT��0H_8���=n#F�NN0%��
D�x�ey�~���e%�V�T��;����tk�2����-��i��IhǣT5�7ۘ ���8Ul�4��؍-�é#8��Z㚄x���<.��C�S,�	�Y�[�r���X�W��I�9^�7 2�v�=�j�oθ\��w �s���򄋠z���$���`S���hIZ��}&�����'�i:�	_;�p�p�o��~�wQW R��}�[{���?��1��2B��Oq�&���PIk���ٛ� h+�9Yp��]m��{byΑJ��O1�c��ʼ�� ��w�VF��Ei�&��{�#���4�Qq�"uO�x*􅍾NG.�\��<��IR������*}_U��  �f���=/�N|�lF<3���O�Z,����s|���q���`nC��`EoU���C���I����P5X�/��K��6h��nhn�_�f����H}�ciO�����aCe���aM	E�Hk���l-	����"�ᾡ�-t�O�fc��Bc?�Y1�s���9����V����)T^b� �UVd�pS�o���ߘ��%����ZT�����qF>����6������-הS$�NIrق4�q�5��D^�6��B�R+��/��G���	�}u���r���X�P���V�C�� K��È�x'5.�KN]�F��_o���C�ɪ�<��SgڃT�X�&bY�n� /?�>�97�d>�ڶ9s�䌗/O3��&74�K�J��'�q uf�6�CO�I&NF��o�3d_/��E"��wxde��t'^�T�nD��&�^����|}���åo��W��_��1���Mf�z�y���ըX���$7E��������%^�i����I2C�>��04�2V���wa;� A$'#pA�1�%�n�%cz���...�t��<����x\���1�5/8vr���E�92>�t���.��y�~�{�,��)LO`�����JLT�ZKH�㱾�<v���!�J܀a��(x3w%��kz �ziZ��Z�u��s�B�JC��z��_bq]�3��=�5!$�(�;��#tx�z�n�q�D5�ʝ�J�#����>�/l��������$-kT�L�@Ña���)LhAQ��=x������|S�x�ɖ�%��)?~���{��A����T-�m�Y#y���$ӗk���ǍwD�8�Ŧ�	�	�j����<<�+�RV�&�ȒZ|�}z�fů��N��fa#��i�o�o��xab��z<ӌӹ|���W.z��l���Uq���к�!M0����	tyC�v���ZL�yo']�]?����2.�|�R��&7�V�����"�q=;�K������zy[˂��o����|�G��yǇ@r�1	���1�)�5��9
�� J��?��T���v�9�$�mNw����l�+Ýֻ��p"�)����0>��Q����a��qL��/��g(���y*H�(6��0d�>5
B��?�
u}%���i�a{���{0O��X�t$�R�P�|��;�m����ڕILO���Ui?}��H�tR��\�B�,Vc�+m0 �f�}���~�"c�&�M��a�\��8��t���\��.v�ޖ�Tvq'�ơ
n��8zv�w� t@;6�cO�p:v�l.�A�̼ݫ�|2�VL|�[Q��ή�<"�@�����P=�s�V�"�)����b֭���s-��:i	�2��.e�|��E��"W��̂i֯�׾��hy&��/�	h�2�U�>�X���d�z����a����XR���֘�,���;^���\��m!�WF���ޘ	�
���%q%�0r��tGm�
�V
�en8ޞ������o�J49�M���=�����-rl��k�U���<�	w:V8O�/�:ױKtq){��B.��_h	�s��܌�;^>�H�XM�	�o��IHS�)�4�M�'ϋ�U�{۳���ȃ	���'��, �=Ó���_�ZѺ�r�@R*:�"��K����Z����pX�ŏ�Z����؋�D��ߦ��2�ΔM�AьdC��m�]�vVl`�YMNw�I��z��P����dE0�}\��[��~>�Yz���$�ůӞ��{"<�ə)Ӆ�K��#~����^"DF�����7�+h��2�뭻�,k��wƟ��
����5�ϔ*�*���s�"�Z���X��l�ӑ�so�"PCv#�3�D����s�d�Ulr]���㿤)�7��N6�%YYOߜSIYvcv*V~(i�}��h��6~L9�M>q��9��b��G��4�>����3�)7��m���a�e��=^S�G������ix�qL=h�L�wN�8 y���i���e�
<�K-��K�lpn� ƯQHR���ML��8E|b�*a7�{݇�Gc)Q�	�ņ����$Q�9�09\ ٵZ\x}Cj�z�.6����ؤ>S��:|1f�����k���3*&��I��	�8}���7��ٰxSs�2�2���C�L��H�wwףb���0+#�Z�ۧ9a��+Z����o"��5�5*�"b������f=�B���~�F|{����UaF��[�)Ά����6�Ձ^��?�Y�?�oܖ��W�2��M~F��ZZ��a�e��ɝ%U�Id�x���~�"z�A��<�I�S��3mi?QFcNZ��E;2P��Y���j��JC�����f�)V!�O�Y����Xy�������N�i���$/}ל���l����7�댩���][�1!�y����Sߪ �03nlҜ1�6���09�V�L
xX��o�=�{\�����ڈd���s=r2d ;��q�Q$�y\n,�GS1�����S�F}�(�l�qT�ʗ����Q ��2�Z+��y�`MH	n�"ۙ�`K�O/�����8o���\�����S�V�/��{�U����.r�T�	9&�5�D�¯�݊'��[�D��
���j��>�IHX!���lS����5��L�8X��c�B�F���6���
��9wJ��=$ZDFX� 2�:����!�sW�m�9�o3>"���o�=���	�	Rm�5�Bu���"V!�G�ˬڡQa�T�B.���l�Ge�aɬC�P0��XF�o�ҩ�۫��q��L�۠�r�-��wQv�;�2���s(U���)��� A�y5�����p3�5Lڛ��\�~�c-mTB$�Z_@���p���p�����}�-������|F�jG���%�"�%���>��췦
�Z�g�=P^�LFu6j�Q��r���)��/� �3��U��G��XR_(���B.��ٕ��$2����<U��V��j��	ҭР�N�kl��}��5JF����ųU���0U&	�u��TǀQW��Ӥ8�=�d��Fנ�����ki	�mM��*AZ{�)�������e�r�LC��������Nny���	=����ņ��4_���Z]���dZ�����따ߖ+׋Y����PQU����<H-�+Ź�ǰ��ɻ�o�Z���ex[����������֪2��5 �/��SV�����{Ǒ*���)��pSJ"�xZ�٦<��6}�}�w�^
u�c�O���a��:>]fn�����A.ۨĦ�Q���ve"�םS���J�T����N2��dʹo�r ����5�b�I��	cT�!5�����3%UV����s�i\�\��:$�4�=iP1L����ã3,cEĲ1#"�ɳ����j�쥢�q�Q�}	�v,0���X�F��+������â�����@O�f���k�Q�2M�h&7]_� �O�k!Lq^���ĥzM�t� �����O�~0�Iʹ�ג\!����;>3C�A�Р�$r>�_'���U=���4����*��AU'o\�\)�`>�v8�U'�C{�=I�M˶�k�i��?��x!�O��F��,���Ϗ���L�&�����➢�9jUj��D!n�{�#��)?�;���rΗ��}���[q�*_n4��E�ˡ����{�����OTo ]�Tw<EK������!��I�Ï���U��w�E&`����U��/@�Nï.��n����5��!�&H����t{㑼�osX~k�c���9r�#���TF=L�A���O]�5����*�/Q��7ʈYŇܯp��0�B�����_�s�^k�J�+��%��w�tEʄG��=���+;�r�	l���F`������ve�Ʈ����{���梚=�-�r)�RLO6��2�?w�Cdh��e�-M���[�N�  �͵�P7��5*j����P�����<|w��."�T�?!�
��[�KBnB>��N3�"�D���(��_�S��~��y��8<�Պ�?���!�h"X1z�; ���f�\�TuEX=Ó5pzuGw!�N�$��]ɤZ����0��'km�!��Bm���O ���L��� 鎺���.��x-�u��%4忹(
C�.L�P��5�hJʓ��� ���a�F�Dݦ����!���,��:��_��v1��+���,_H��%��-�{#/�����I1:=���[�N������T����jkx�}�a����" k�r�u���/��/�"�G\���L7.���\O���
{���R3�jE6쳶}���S�c_�c�6��L$Iח�C�ܮU/�j&�x]qk�SH#6Rp��`��x&<�,���AN�I&���MM��V#Ҁ��v姱^����ɲ��
e�_�h�A�,`���b1���A��k��,���4��{�5� �	+ߞ��v�=ĜkhepY�>���^�ا�G0�P���/ז&���?�qŜL�0T�B�7�iv�9��k�����6��߾rח�:*\�,�,��
jh�xݦ�����9 ���d��Ŀ�H����Y�耓x2�&�ʅa�mKn�L��ϗrA�Qb�}5����ߦJ�r������8�W���U�w�ϯO�4��$��=���{�u�
hF.�ɜ��_�U�L�Z,2��g0�Oא�ڈ��tE�p��ڈ�����*|Ο�jS�םS(�����A;$[<��_ s���i��^���05*wl>�u��Ĕ�<����n�,����@�lb6n/E���ma'�m ���`�u�飽D�����kk�I�:����V1K�(�c�
�RH="�d���1��M�����Ot���]�⣵��Q}��I�=���-�lפZ_�0)��Sc����8���Iv6gG�G\v[�3���� �Tq>���x���c��Eg����7�U�dPҼ�'2>e�I��Ti�=��j��?O�"�H�OK��p(t����iD��D���΂N8�C����/{α�Po;
Yv�[eķ�a��������Bk�� !��0h �����sx��m�0�0c�y�c�fO���|�0�]�)>ZJtW?1�؟-O��wux<ҟ#���&E��P~��.?��2�Y.�U(yc�\.�����R<5�Σ������Q���s��xD_�0�T���Ym`�OE������fuy���}L��WF!���vN�q^��U�ׁ��%�$s��>xj��18��2� &��h�u�	����ohk���:l7ЯE(��̒�l�L�c��n����	T����'�������dS0s�Q�B@nr��s
�Ew��05�,�v���Gt2os스FИ�� K\���`kC��b�eP)+S��"�Hҝ'ͫS�Ȏ�<�%�h�y�Qn�ާ2��C�:�A�q�R�~��L�ƭ�4�<2���l׳�'���_A��2��XL�ɲ/�h�?U4uze�f�˶��6��v�q�y�<�r��q��ј@Bu2����_+���3ʤ���g䌳���t�Wj�|���&N83S����އ��DJ�W�sJG��\,��U���o�")�@2�~yU�K���ޑ�g $>��q�q8M/��d#q�u^c2�kS�3xX���"0h�(���343�(��J��
Wmܢ^zc��|�]�b�)Կ�+��%D�f��D�;�(����jY*��gm�,�[�U���m7�6|5��<]�5�]�ȷ}�������~�െ]JX���ր.:��f5o�F\�f�&�m,U^����f�gGނ�n<N��"5��R��D�W��19���U�#f�h�,.^!l	�p�Y*��Q~���S��X��4g�\���&x~7��o�ᵨ5��QcHuO���w_O@/���Y��� 9~szL�"ߞ#��L�~}��#c~L�X�/eז%2b�&w�&yM��7^��̘s��/{[:gE�io�O�#k$Zb��:Z<��}��	-�r�U�z�ח�|w�����p0�V^�IL=�rJ����?��ͱ��]g�I���&��%$���D���@��Z��fK�|�)	��a��`�O�0�`�t\�CGs�q$�����x����-=�m�}-}qY�~�^G�=Z�Z�]q�<.J	�j$"��\-?H� 2L`���p�����'ہ�=w���
@%�*�G��0���y�³�$ΰq�ּm���wB�����כ��醩M�_ۙ�=QG��� 0�lP�@�%�m>s�u���'��<� M(�?{n~6ߵ.�]��0_���aT�҇�_-R�ɾ�Fλ��l?�¨Fd^�;�uTZ'=��,����E�S����1<�o�D�������F7X�N�	k%kuz�!�^W�=�P�S��ϗO��(�2��� {}Y3:s�M����8��q��*��/��y�>�f����y�)��2��|yvq�)kJ?>��
���˹�ʿ-N=��餋|n7ļkH��u(�V(�{�α�.2�a�ٳ��Tf)ǽc ���ǖ�G�RdD��n}���^��{R鱧/@9�5�-x��[ A�4���(hC�Cb��D�<1�Gmɐ���)�T�����5*!�rci�������m���**�9�E����b���0B��n關��z7�Q��*KY��i'�s�]��!
#S�v��#������8�.��B�8]�h�MR����*���0���.r�ܔCAqz�Z���z��g�,[wY|g�(�U_��* dܸ���>���mcy.%V��+����?s���)�Ғ����0}��G��yO���E��\3V��zҦVZ7��f���V��}2����
��������u��.�
���HX�
��F<�t��|���BIm$6�t�"�?��Ms�:������W�G�3r��14��(g�kH�+��Wk^�*l��?�{��3��X���n�ct�y�ON>�O��EO��R�;Ғna!Mǐɍs���c1
��{JI�G���k�K�I���"�����~?Q�5���J�����e��'.ߤ��i�O��� �?92� ]����}���_�Sx]��0�#Ht����П��`���϶�^�5��[xL<i�yj)cu�p�L���݈j0]���j;$�����w�?(��|�]aSl�ȣ�Ba7���ԧ'���3��`'���V�j�Y��c�*y"��qw3��+�������ޮBA��ŅBt_i9hF3g�תʄ�	%_I�?�����<,���[ە�0ბ %�E^l&�}�ph�J���2�YG������^�<ˣeL&R�_k�o���c9��vC���f��x���LBZ;���D<7�J�ߏT[�6�Gm���8T��T�����R(�h��G�7><,����䄻�ў�mg?�@%n�4�zL�Ov���D.v%�~�4og�w��6�.2G�p�B��uS����1�T;��������ӜY�ڸ��5�X��Q
��^�d�)���x7n�K����(�Бi̬�/����L�m��yBɍt� ��&�� �;���d�%�VӚDq���O�Ϣ�}�ISk��K�JH>�]B��U-��!��٭�&>�1O�Q���.�����CC	��C�	X��D�f�EG��� B��87z�V��W�D��x��9p�a��rӇ�2�9N����6�����Oψ����|`r?�x���+C
T�S3}d�{�����3�8ZZ&?s�q��"��u���{���g9OTym񘛸����2�I@65,��^��[R�]n���Z�'��;��u���b��qد�����8� �
�aL��L��g��̱�o����{�����[�<U�"�B���/l����	}��_Iy\�?�{�;_�����--A�Z�u����yb�m��0M\ ��p�^���	�4�vDv�{Sڲ�n�xLs�8`�qS�UR����T��Q��̟�U,h�7�Θ�̹[O?�Z�Z��3(�"fwoDm�����xǡ�m�h����X�a�8OS�	?�����K'���;�|t{�gp�e���c�uXW���)��l�z��p����I�}\�1�=k�uʤ�04���m��%�
�*u��1q+UE�s�'p�^Wn=�������`/��fEl���xuE_��,E��w�`�4n�2_�4g�>���P�ڥDg��i��R]�*nT����o"+�u�f����H��@��ل�Z���F��v5�v�H���1sB�Q�1��V}s��Қ�׵㭹z5^����\�#k��e���ȩ@��}8�f�I�"fF���������+�[�n_�;},�`�����KEj�O 4z�*<���X�A���झ�ݝ{��ÂO ��F�KaOY>3���>��5����QBb���AQj^����ޣn����l�z����L`N;��U�KĢ�k�
���Ku��RT�g�)͏�!��i޾�sT�O'��#��G#����i
O��7�@5�N[�)�v���=���On5{n&N��R�}Pי��=&A�7�ϭ���#�H�|�f�N�I&@�T�����
7��D���fĴ�_)G���w���������jrk����9r�RP�IWQ�HD�(�!���L�  ]�=jh�A�H-!t1�B�y8缳������o֚�<���.�u������PQ�
7g��D�������B�_g��j[��qB���!�5y�/�g�U�P�˃��[4�����Y����ṯ��F�X3D�����n��e*V��l���!�<<'C}�fg%� ����� p� �P��^�B)j�?��\��\������|����n�{чK�Ȑ����x�Jն*$������rG��̢z�8�Qmk�{�9vj�sY��k�Վ}����o��U�Ϲ`1/��<�Fv�W�cY���ܹ�������>~���e<W�~�`�^=�U=�W�D�M�;3���*� �x��K_��C�4������uӧ(�6o�zf29�6֎膿�� �9��M�z`�!#�9�������}B՚��,C���Q���c��)|c���}ҫ�g��U�Q�9^C]/R�U�������s�ŎUx��r���pG�A�������w��ß�~g��vLTF�y���5²!��-6�b���1���x�&p\�I�{�^�_x�?��t돤�҅H��H��~�wl�|vU>�9�k���xB����e�'4<���7vҵ|3ɸs_���w|��W�#�UM�l��Jl��Q�	��wi��x�u?�L<Z���6�'���"�Lx�D��Q�`KˇO�!,�X�>h}_��LC�j�ّ�֑Y�$(��!���t�"*��_��SPyֹ3���f�.���;əp@LWfݪ��0p7�u��撥�Wf�Y�aN��X�]܀V�F�4,9�?�
�.�d{����&����i���Q�M�U܄M ���Ym>�W?����9�Ӵ�k]��u�7�J�0��"'~$X��t��K�V}�JR���]b�2�3��Jd:g���r���k�d]��Ĕ�ڎ�wͽ�k��n@��b_���w �W��×1 p������M�������GL� ����t@-���{j|!���e�\�8�48�����Քj�<�/,Y�K��r�̖tz$�H4���L�����M�+`"�����S;�4����ؤ���4٩8�k�&����ڈ`����@6���3����s��[WDl�ȝ3l���t�8�o&��Lt��Pa羥Z˕A�H��N:u���\ bS����v�͎�>����ۏr�U2��R%o���d�b��czS�U�ě1�L����b�r*u���c� ��%�q�!
�٬AGB4YU�t�4�RZMw�j	ݻ�"G?��2|�����Z��XblǺܝ|���I�-�9������8��ae���m�^D�=�q�a9{�/'x$6t��5��Лte5\���o�!g�[ف����Gt�ֵ¯0�g�h�o���ܙ1�;[���{!9a��y7��+E�/�eG��, [U�V6y&�J�Mc�eOՐ}̋��Y!2GBE��^&�]u�m�a�7 �/��]�5��8���m�4�� ���������e￤���a���c)�Y	
�O��du��S �΍KI�uA)�y�P���^��S�VqZ���l[�&�:�j��T�,�$���5IH���9p���g��me�r�]aW�y���Qq�͝R�U/��T��|_���q��\?�'y�VZTl�,)*q���.�����yK0F�����`4�I�@~�s<�
���2Z���Um���0!ſ8����!Yo_��"��`OQ��D��g��h��.�4R.1~�t�ė1V��nݕP}�9z��)xI'�"GĨ��"h5��Ǩ@�[�z��$�d5`�Ĝ~��ͫX����ʇ١�������S�A��6��&��}�}z��A8ܣ�D1˛����q� �M�S�ZFV��ؾ��%�b%��6:+7��`�o��Z �	�.�y�U!~��D�ݵz_�������7�8�Q�����]m�ryq�e���gu+�	 (d\�F��u������K�����ɵD�m�S�6y$���I�Y����P�6`��}ӷ�k=�c����]�/|���Td*�"8�}�I���*/��,[�"l�槅3����o�",c��#m(��l0��(ON��C5���ww-�}�{�ez{(��wX.1���	\��LXU""�#�oʇ��x���b����W> �/wa+r�K�4b�ןD�m��:J���MP�m������7�Gه��N��T��#e=C���Z)��&_4jX/�Y��3�l�z��r����V��E?�~&���y-R
������)�q�
�0*`j~��/�q��LZ����&4Mp&��gi�n��!M���/�"�l�[̺2�ݷc�)?��P+�q����h�S������j&�o��{l��ec:,��ߔX�����AK�6���rG[�?Lq^P@��m�Ȅ��ލlEo�fb޸�)hi��ƪ�7�ݚ��gn�Z) yHk�_������X�E��_���s{ a_%�T`׳W5?Z}.�C;xD�x����^��ʀ���8�!�CV=~j��EJ�]Aw;����~�]�F�����>�vq�1� HEHY%V5�z�P혡�Y�|�^}?PӍ5ISpU���ѵ�6E_j]��͚���-
�Pu�u=1�3�m@Ц�WWn-Mx|��"�7_��y��ј�DU6���N�Ho�m�����q�>�Y�c�6�ޒ�t���w��4�1�K��f��zӸ���@˴�۩2�?��@im�Sj����Yr��c�D��T�by8�(��?��q�:�!�˾��42��TSҔ8�cI{�P0k����_� �M�H�
�g7l%Q��jw��:Y[�.<%�j��"kSd,%�6D\F��S��h���e5�}k	���3�i����S��HA����fϰ9àt�y㣭��"�89���:kn_;)k�s�<�紷O�(nbV!�̖�*�E�"� *����i�6O���o��D��4H<�.N�޹��ؠ.��e�N˵�F1J�1O.�_�U& 2)Fc��(�бґ�1 ��3��fF���$���d�������gJl �t�h�/ݴ�O�,sPvz�'/{�������U�ݠ�H��A8��P���8���)K�{��i8i��Ȃ��6s�AZ�u�#X�7����J-Q�Ɨ{U~���v'!z�n ����I���*B�i� y _�&)�G��/U��cs}�S�∴o4�5	,�R�\!}Z ��^��u�����h�I��X������h��4��H���gW�on'9�GHH�+gv�"S��J�{��l?�YM]�]	��&ܱ����������#�:�r���:�e��R�P*�zU���5��OV�g���jZ] ��F[�rFv�7�,���-��KM����%��5 �
���K~_��ji��F��F�q�jW~�c��G#r�q�g��%�e��A������`�i�
�s�]�`X�t~������ss� �q')�*�j�~z�,%%S%��^5���.5�+�`}+����V�~�G��vXJ����L�$2<)��k�>�t�2�����ͥ\i�#4|z�^<R�8*�n��l��]�U�1,�l���Q�̠{Òr�Gkבw���u�
a��b����R4��̪�.��8�*�h�7���L����q@���G>��ןt�a�W���9�'�oC�E{F	Hx2��:���_���RH�rW�j����Z���O>V�\
�q��_�=�.x��*{=?��0����[W��5�9���H:N�BR�1�ɪ�j�cb�+�y A��t�9���U
 0Y?Z��h���m� o_���� қkv�����GK��1�ha�3Ո�jK�������u]�e��s���y�t��Lx��(���ˏ�,D�rܪ,O'?>�si �3UE5�&���~G8��a5��4�ޠG�Gq�:���˶V՜��Դ�G�����'S����X�����2`T��^6��~���=qK;}���Yg�u���3T-UM+��9h��|e����n���A���|-��m�;�Í�����9��l�M�����x��ԟF�h�r�M��/�p!�19?�^)*��b?�(.
8{����U���<5|+��x���덵�I�VX��@����dSz�����ኀx���A�j1�z. (`�>X~_E>e5cI$֋b]�b9MՑD��n9l>��� �t��AQ���r�W��	��o��.%�k���]�m��ț��Q$��������<����w�e]|K�Ҋ&e�՟�^}}���5�,F�rUHVm6>g�8�ԑ �t_�U�[�H��5|��6F�5�I�p@�y�/�ʗ0��G����8G��n6/U�FW���S�&(	��1 �YTX��L�ϝ7� ����1n�Yt�A����#f�p.q���;!��AiOȀ��ٷ>�,�5�s�5WxT�Z+?�=�B2�R��:�؝)u��o�}�)�;��z�-�/caN�]��� ��(a��]�Q7��5�%�2�8|��Qz���<�SvV%�:Xp/wk^�4�XwE[��!5�O�>}23��,�.�;����/��!���\o��hm`�Q��)����uN�u,�d�GެdH���|T񷃇7�`A.�������4)@�}�ʣ���G	�K	a�ϼ��r�9�8-*
����{Du9~2�{����L8��}�H
>?��t�ݣ?���������C�$1;��t�cS��@��puiO��B,�f���D��YP�-�aIY��xJ�5)^.S6�Z�8�S��;��^;��t"�<�M]��"Fȗ@��A+mΨ�_��9��5z+}�����˾�c/��:�w��D�e��r��-�䉷���{8@�}�ٓ�fT�LͭbZA9���	s-�Vl@���I3:Py�����w���Uu�HGX:��ݤD�T���j�@��k�Ҧ�ܠ����Z���C�9�vD�Ļ�S�=8W|����<��J�p������gN������~���M�^4
Z��j�4J4Xo�����f�7F��߭�;�8������	p��&ݪ�Uό��Z ?-��[�i2�=0�d����#:@:L`������&iӤ�O"�nk�$��+�gm;����0(\�I	[{;����2L�9�b0b��<3wm�Xm��	���8��� `��1���8���z���F��i�MjYH5�G��j=��J�7",����-,�ļ�ӌji�%�,!n��XTc����F��ru� zg�*Lb�#Ζ:+��!g�W3%bVu{�T/�d�/:�S���Y�E@��
�.4�����mJ�iI�Y� f��
^��+�6ؖх֛�b��]Z���$�(��n���(���ͫ^nZ���\�G���=��ńU|�l�{�`յ�}�"��̞�gV�8�{�k/�8��6�02���y-�$�'�a�V|.#5��֥�[u�q�%�FP��d�^�y��q�;�Q�0��?&��D_
8��'~��Z#qc!f`|U��&rasƀ��BC��K�'�ۚ��f��N�Y���4�Go��7��Ü�k�o����p@w	���6��ix�nwF�i�ـ�Z ��Htf�>�I����ގʻb%�����
��9�%�#����ez��I�u򨆋]��}  iK��6q�y�4R�Y[���հ�<�����1l`���8�-��!v���I�����CG�v�҈\]���|-��f��am����o�B��
��]��,˻w�W��՚���M�r7(4����-	Q�_>ӡֹ����GNq��;�T�����w�����T�;1�!��Fak���4��L4��U��m�H:���.b?���-��fK�3<{sĮ)�>p���^��'.j��xwb���
��k�á\�i��[�
�|
u��qaW�H�B��q�t�m��Etx�pdk��ڼ�X�h^�u��	��#�x����QK|��J]t}Q�l��a���=�^w�_����J����C*;� ��[�3>d�k���p:�c�W�E�Q��ǋ^z9&���T�nHF�u$�(�)xk����ҫ��������UO��pY�.�����o0��%C��{+�p��n�TV���7��l�Í!?1�$�׎�ey>T�S&�7Y�>�%o_&_d�K=�z��S��Q�y>$f���kw�9��}41�A"G#�1����:�4J��z��烏��������gyM��� ���8'�l�r���e��<�N�>?FI��2��
��/|3<3����TZ���p�Ƞ��B�2"�Mػ�X�3�љ��Y�h�?'ez�kpa��� �bgA+Ymj=�6��^=�O ����.�k�??z��F�-���0SY[�jg�}��ѥ�gU�����&�P�+�~�Z�Dv@��=���K}Pc�B�����Ŗ��{mˤ���O�7h�	���f7�3 |���V�(�O��%���˛N���=�����~!�B>�)�,����4�!-d-�rc3�Aߥ���)��r���_Ы��Xg�}p�˷W�EFE!�_�����<`��^#PVu8�<��T������i��3�4�9���Zqŋ���L�9�vHi�!Þ���Ĳ	�<^jC�4
�9S���Ɇ`�����7���@�߿�����j׌�CCr��w��B�q���+�}�Ϻ2��<	,��)[�⡲Gk����k��s�XD��J��X�\���P��"�w��k��pD�/�uE����?TR�ȇ�߷�{~��p�	8`N��� �o�b�ƍ����u���]�jG�z��v@P�][�~���`�B����%v�`��+�x����t^5�k{c�ng�e��k�$��4V[���K��I.o�<�	���(J���.�/�IA�b�΍��e��,޲��t��Q["��\��?�b�'�{��4JD:���&}�vr/�V$��l�i��4/����OZ���}q�k�l��[2�	-�%$�1�w�6`���uo��
��g�q�- ��ȁu�KM�үF�k7���3Gk���O�MT�h�p+��?���?Q�D-ts9�5�'v$�s�;�dἥ��>uc��߄�G�H����O��q��Y��.v$z17�'���E�/Yug!���
f�`i?���bop��[��9"Uoc�GWp���}��ڢ6,�Pw���ٵ3�(�.~#���݈/�o��V�����2l=ve��I���x�4+���9�M�?}�ґMoZj��|�Y���+�� -�Z��n@ ?���q�^oC�b9VUzf��\������������B =t����b�S~Z�yqFƓy�������ϑu���O�:�O�Q&Q�<~}�?4ĩwڄ�zo�/_��O��|ރGm���͑�ʏ�C,�����ٛ��܉�^��ޠ��g/]zP� � �㠂���_�;Q퉒R�ݮ���R�	{��Kμ9�q[�Yx[�/�W�����Aq���+�o��4��;5}��222	�����յIxg������6K��GQ��q�3M=ٓkfY��^m��\�x��F�\���䵽y%��J����,Ǳ�����,Q6ɵ>��E��<���E1���|&�p"���|22WE�8�8�ۤ޲^y�x��K�|�m�t��Ƃ:3CR�<����������"���JC�P��pxc��aj�<{d�*���#��0*�s(8��u��y:M� I���mK��=o*�Z ���0��v����&1�m��6
��K�4�������
D�y�T2���n6?��Og���;h���\�����%�0�leصk�g�|ʎC q38,W�<�y��]�~���:'{�pE& J�� wB$=��(�������)vw�g�̌U ��^�2�+q8q� j��G�o��c���W]ʱ��gv!M��;��W�(�x��Z�L94����y�Ov�E9���'�׋���w݇��J�����B����A�-X� ��iɑJ�֝X���c�nk1;�-]����㋡	n��B���E_/�!��Ԟn�Ihf�M.	 � �>(�ݕHP<Lq��͐���7|c�s���"�����U�o]�^���$� ���3=n5�L�`��#��+�oTX���E�%)��P4NV�%{[.�o�=��'�6�oE��R#vC��C"�\���0JS�8�K���
�O��f�y`Hy�����^��&n�g�_癮��IՋ��y�(.z��\6*���Lz	��=��m�2<@&�9? ���51�i�ݔ�k�6�1��Z '�脮�M���.�<��i���47�a[���5�<�C�9حI�ەh�3�� �� +9C ��۫=Q�0{?���&��3I�V��[��#8��g�@6��*6�Z�'2Zqۋ��	11`�}��i/?m�^���Gv�̍���{����0f�U��-���f*:�(�Hr,ȇ��ùb�,��L�P9p��Rpu�/"���L\�έ۷ۜ;'_�@o�@��{��fl$/"E�t��~�^7��*`#�J
_���Ͼ��P�G�e�l.D/�~I��މ���<Wp��M���I��eO2,�ee":��ζ�v"$w��J8c��!K��Ke�!��?	�g���E�Ԭ�@�>��w�R�su��)�פ��\��&%K���~�[��+KA���l o:���k^ `�,:�(�JP��`��{�X�t�w�9�7G:��(AZ��l���[kY>Һ�Uqq�1%D�����_�����i���
�.C���׼���Y�&W��B�:|� A�X�4m�:us:=pqC�8+G�^��t�y�s�7F5������m@9o���۹g�z~�kgkx�Yu�ʽ�ۍ7Ϭ�I){�Q\5��r�ح�}���4SM�^���;�e����E���fi���f8�z?�	��=Z�D<z���YJ�s�����໒,@��7/��UD���+ N�{V�]��r����/}Ț�Id#��?o�ޓ�s]��O�u��V��:���@�*��S��	�,=��f�G"����p�p���˃�X���"����=EM��~�/C��~8J�����Fk�u3�#��x�3Tl�DP�w���"ӅW��s��pĭ�ij�^5��%b?�/��1v��C	)0�ƒ3|[ůP���#�&��.aC;���;��s�k�3��m[#PƐ�Ə��UٯV�>�ǘ?�d���/̣�2�u���1��[^'�>����`|��^��-���v5Z�k>�3��>�����'&�2�b5g���3��c�)m�Dq� ��W�ϫ�kl|���6��-С^֍��[w
kIA��|�`1R't�#8z���H>�#��o�Z3vL�����7�BXz5�1���ꍲ|��hH��o��i
P/��wN��������3cf�����T�o���
�?۬�5?�t�)V�1*d->��
�g����z?:�59!��N�>�{�k�۟o�`�O*�|:�
@>���K���_�������/RJ(���h����@.����ɡ��6V���G[���(P�����t ���^����h�|�������e�/�5��Ĝ��*{]����/�돏,p��c�N����BZ�S�k����'vDT�Xy~�I*��v�晀@;�H�MR�t}U��'&"-L#�����(!} ,vy�q���Q� �q��h��g�X�N�ȉ�j�C_��n����Z���*e�G����g_���O�\Їz��>P
�R�Kw���|D��ˣ�j&@L���V��;�4� �� �+^|�J��+��$9KGwA�F[�����H�y��m]�1M:v�p4��zg���̗6���@�㒳{ ��*^�H�,;hr����7톮�?9��!`�nI��<��sl0B�CL��̴�2�xDO��'(H��=�A�۫�dZCD�]�ؕ0��3!����N ��
��9�d^���`�� !ngJ�㈊��<� ��ѝ�A����t��F=�k�I;Ӣ*�&��ՅL�D�ѫTi�<[vo�I�w�lk\<����}4�b%� B�ϢA>�}>]>��ي໨਌z`d�f)"0����͹g-���I�:_�9=
��}���^kF%}��~�E}����CXp�п'5�@��\�(<k�n�D(h��<F����a���E�
	���|N趨%�8���& :{�A��G�o��FN���BYYd�^,>ܑL�j�w-� �VV�uacy��|/Lb���3!�95��4Z���>�������,o �kK�8���$�vS��a�9<U�����ĉ#&�����*�o���TE�QU���(��{�pGV�돇bm�*,%wg�ʛϚ�������M�]�"��O3�{�TUZ�����i��n_"�֭�a��$px8�O��]-�.���3��C���\�N	�����w�}(��^������x���&=��5Bp4<��ic�!a�#�]S�Z*4t�L�Ƭ+���kJ�xf��­�@��Y7�o�����iQHb�~�%t�M&�Ĉt&�܁�LD�}��>Nm�p���ަ�����Z@�I\���׬r��ol�>�l5|�_�D����^�|>���Ϥ��P�K6:<�>XTF�ȶ��蠖i��W�M��r%l�����]� |�wV�߈����Wb?��35�&���.�7�7n�~�S���de���
��_��If��i?z�p�R��~1h}?��T�`���TO.ع=������W<Zh?d�7��s�)�����k+������dfߛDf���d�h�8��
�zZ����u7i1���/�F��c��v;�Ҟ�b�/k� g���[��xK���b��L$���MwX�1�#>��ZZ*��cb	%�'v�)l/ ������B�\�� 4���i�0KÖ�K���V=9*>��ox��6C�.�$-F��E�h>�M֚�%����	��#=ާ�F����P����{&��-:RcDSρ䕼Z�K���XK�`.�n{TU�w���p��^Auo�eCC��5�,b-�q�?GGN�̴��:�n�~���� /�Z���p7����'��8R����(Bt�=��m:��-��8G�(c~��ΧP��+3Ϻ�'�1.���ބ�'��=d4���!��sTܶ�q@���NsJ�/ο��g^.������(� �49pQ�>l@Eb�n�;�O�GT�bw�n��2VѸ�ʤ�K݅��큄=�{�p�����.aъV���d�`�4��0 �j������N�Z��~�pʃ;иZ�nv>����_��' � s�:����� ��y99m�=n�1'�"5S�ܓ��k,��k�h�������}t=Gg5����\�ݔH�}��ڥ���C�Ҕ��*�5w[J�~��n�����v�^����S=�0�'�����dA�Yh���^�i�� ��M�2�M�隋�y��g����U��l+��V�$v�^���*b��5�~�Z�7̻��a��~�ޅ�|X�i�j�>3�����Ȓ�冧{r��ε�&��#$�`�A��s𨜐�!H�T:�uRv�RnU�LPS�]�"�=�PqH�Q�,�Š�7p�M�:�W*\���P #o���Ѱsd�o�!����N^��h������Oȇy�/4���Qe�qp�(��Vo:�d���oH���&[�����U������W���c�LU��Fm�혟8=��(��;o�5�	j2�ʩ�{1��~{)�l6g~E*���C�������K�9u����f�&��mmU׀��{F3�n�"M�$vVZ��! ����=�|+�n�O��Ζ*-�U`���`����j%�$]O�{��r�R�$m�EORC����|$p�Jw�����ɞ*������ZC��D���m�Js�֗��Nm�j�>����äT�	H���Bp$S|��+�VZ�Qx�BI4�ɶ�AHX���*�^�7Q%O�Ы��͙<y6���*����i�յ:f��^<����z��0a���P�īU@;��O]���ҍ����������M;_��-���s �؝�>�'��U�=a�S!)��Dr�`Ee��c��qg��!�ى�x#}��E�#�Q�g��:��&�w�>/�}���W r�U�����s���>F����w��O�m[��]%|����k�A5>R$7dmm5��o��� �`d�ut:1p�JNM'��c;x4��1n�6s����vG�ٯ��9�d4Pw����಍�9���uO=��+�.���?�?�&��z��&�Sw������">qh�}RRd]�IsJ�e�*�PQ�k����e����Q��ܑ�ͫ��嶽u��/N4�Y�f>I����]�'��3FsF�4([M�އY΋�����ʂz�rrڑKkkT�:%Q�;^ȫ�d����؆��ѣ�a�U�l�O�8:��𶢚��S���r�5�Н`K�p�Z\�NE�=��PG��w�D�2�I�nfb���vp����p43���Zެ����&���oM�Y�v?^����d`��h�g���/���(U�nU#�:�O�[�+8al�&�����׫�M8�������ƞ��/T�m�� b�]���'��o;Ѷ�	���-Z��D���S+e#_><�t���u¢J�6#/p�zV(8Y7+~�oS4��}��]Vu�3�d̵)�VTTx���v�������j:��Od�V�;ۛ��!��n Q��.f�uߓ���}��}��Ķm��5Bz:��̲��L����rh�!�:����"R�O9E8\��t$2�~ Ҹ2��Ϳn	���ZG��7�����b�:rX�G��PJ��!	��;ã�oQ��g�z��]�* �?�&��%L}+y����[�w�D�u(�Rϭ��z;�L/�o|6�`xhb1g�\�|5l��|��}��ݶ6䤼(� $������^����v?M�3��Dv�+��g�����g#��%W<�� PK   O��X+���  D�  /   images/5cebb09a-e86f-4cb2-800e-22da09d26481.png�yTSW7k+u Z�	�5�����dK+�т*�"�2$�!L�
���QF��bŀ"�@ ��IH��D÷Ͻqx�����w��ֳl�9g����>7湴��Dz��EA���k�6�������o��*���>?���=�'|^H�{؇@��A��W{j�<\s�W۳6d׳�c�.*��v������E���/�_K l �~�i�����n?=~�d��y�>����g{�.߱�k?����n��������k=.����yAʶ�S?7/ot�Qi�y�u�̿�]1�����_y�͜�~��z;f��ln��	�	��To��*���w�y{YJ��|���\�wr�k�0�g��2)��@�0��P7`2E��]��Su����\�64��b�BU�c�C�qs7E
{�U����|�
d� d��\�դ<M>��ᖼ# ,��m���/;K�5������k*�pnyv����ßM�GV�m�o����߆�6����m��m�����	�(e֚�ܩ�wW�^d�����RX6�,H$}� �o�h��x���X��p͎�Q���cNKCnBI�q�=qHi�e�{O�1=
x�k��U���m�n�$[G��3(��S����(WX�}�O��	��@p�9r_�6���9m|!�X!?��5>B?k��9���<W{���z��˿`��o�_� �ix�2������{�7��k��{����W��r����BE�z���V���7/��e:�I�ېc��2�?�)N�oL	G

�������/�O����"���<�Ot�"�<��,�z瓂]ǿ�ϡ.K��l�V)�8K>/��i|bH�	��w���*���w\ &�[��F��Ld��4�2��f@O���Ӛ�h^�d�+��K�������	(��S�|M��;) ������F�gAB2/	?��{��8y��v�BX�-���"]CY�����i{�\���D�=��j0���f�/q��!������M�u��>��)I�d��dK�nɁ_����Xދ�9s-0`�R�c8�@@�5����5�/$P�]�ر� �tZ�J�+R*9��|@\��5��v?��>���:��:���$2����Lb�z\G9��~\��.'�ny��!��-�q1Ș|B���_]$���	������|oS X&p�mW�c��~�?���{@�9�(���uX�MH�-�0P
����`����$/�������1��1F ����7r)D�v�s��Z|;�\h�D,1W8���gƚ���8f|��J���W���~!Řn�ŵu<��K|���ޔN�]�.�v-��r��7mrue�'q��L)R��+��¥�����z��ϑ�g҄DM�f*�r�Trܒ"S�+�#�+����ϝ��f!(7@?���9�#�?�}�+�a��כ�+��EL��\��&�I��}����I��]��g\B��Xe������)=PI�Bc��<�p��Kb�DB|~_��[$� �Q��=��g�����I2�uC����,�=0�����霫�3h�����tG��n��!�Y�^�&��~��"}d�}vxf�=<���:�G� 1��3���`�}n�ϴu+/?_��nF�޵��D��x9��k��K�n�i��+�0qa��1�y�8��h5Wb�م$59��C4����.��9��ӀT'ɛ�<�T�/�'6����~�򼚄��)�YT�\�	���)���/(�Ye�� ~��J]��*����-M��3H1�nlش-�{	0�`{7i�$�d陼'��K��R����ԣ�����]�QG��P.N���2��;��/��~%�mRN?f��
���<�WE�s-t 
��v�Q�`��m���4@FfUyrv?�m�))������-�����2.nxJ�Ǟ��߀^OJ���X4F�M 
�m%	maz��k�j���O��� l��fI_6.;�G)E=ΫM���/N���쳰,F�Z �z؅�n��?؁��< ��S���¤�h��Ge l4������,�nY)����i���8���>c�7����x&|Ό~LNߖU\��*��9.�S��(�5����^����@�Wǯ�*�Pq��R��ySL
����oâ�z�T@�� �ǯk�.�)�kD�G�e4o�����o���UT%+?5�DO�/�pƁ4����}��"�sS�b,�B5�/X�ٛ@Gr��!y�6��ē�M8�7�I U��� ��[Z��B+j��t�|�2s��R��I����;v���Eʢ:d��ЙT��ob���l�}/!�0�_P�u�[��gߊ2Fu�܂Y��.�T�����f�>�g�?�nY�������g��Q���D��R}=ax(�^~��?06����G/�v����p}�37���o�����s�"e��X�����z�l��cZ/�)<�u,D�Sܮ�E$ �CWL��U{��� DC/@���PcA3��$Z��{7�(����a�]*'��� ��̛FP	�g�G��S]D#=�
}V��.=�칵oL�\gɤ��Ìl2ܚ��N���i��6@KI��7U�>W��ʷ=�i]����Y�ݓM��[�{���ީ˕�ח�>H�=/@��kg��4�|*πTYU/n2
9��֕��^H����.̥OL��&�I���{����]��Ш��k�y[���X���d*���D؆-.*��}�l�U� ���Q����l�e��e,?��b]D~^60V��4���Ӏa�̟�SB���py1�OT�78���-ߎ�5����Dx~ء�,>@�jeSҼ���������rt*�s�!�[ͧΊ/S�F��x2�A�G9P�GT�� ˞��@���'��F�L�W1�u�p�X��YAR[,��8'�$ 2����0��o�=�
		Z�/�dvWC�O���{���.Y�4w<Yw� �Ke[�v����˝���Y�Lw��^��5oW[����e� 5����a���r�/��Rq/��.!�kV�����#��W7�h����S��k�|�Ю���)V����<+KbP��i�,2t�=7�����,g�r�S�4�՝j؝�&���X{L��^�͝�H�����浺K��,=t����O=��`=�k�i3A��xM�t�y��W��^�����O�gﱦ&��~M�pG�3a��f@3H��qo�[΁���ﾡOm%�Z���53�9o�,E�aXĿ/����Bx�_f��;>�B6����M-'�x(���];��k6*3�y��"�ץպ^��r��r8e:��M��%��G�F��E�Yӯ&گ����/�Uk�_祻����}I��hi���2o��6�^��_7U0���p�<��%�?LD����л����g(������ ~O�./o?r�}��y�3��Z:V	B6��U��3A�u��ʨd�jD���\�Κ����ӓGv��n$�[�l�} Ȉ��H�H�m�O[ó�3MI�n�Y~X�������F�A�	5�h*���U�k*�B+�7�Ŕ�(����YY�ɩL8d*Æ9ߦ}Z0A�O���N�'���r���Y9S��wnC+q�������2�>��N��R�5y{!wK��(��x�Ӏut6�^�d�_&őo;S�M�wQ���}傘ۗ�v��?�����=�2�ϛ�J2A<�#��nV�x�[��� ���]�9�]��z���,�:���Llʖ;��� T��3&�_����^T����2ET��q��N����9}�O$�[��v� �͕�,Q�̶?��܂�Qp.��8��uE�B�%5�X��nb�W��j���MY�"���U?~ j'�rA����p��&�7��,�0�Χ�K�P��sE~�*�ơ��r����ͬ�?�Q�i7��̏��:8�H�2�9/l�(H<����^��#�$;�G�z\���,��t��իޗTV5���^���l���|ϝ1����v3�[�9+�je�ŕAc��hk��R�����'@�h���FM��m�	[�b��`��baW�a=�((��2�or'�T�9�pZ����]X��,+.ˍs@+�{e
V�K�n�J�5(�0��P�$K�Գ4z�����wK��nO,!,�N����k��SE�j_��ƞ����z20�kT�l�3������}�{���R�A/=&n�b}�k���8����f��YŎ��DU�?��n�����䐻~ؘR� �j�[e4�;:�ye$"�C�w(R�3�o��9���{���=��:�6"��x��
k3������Ṗ�ɑ#p���ͫ���?12�^m���'t��2A�f1��Rf�M��h�	�D�:[�����h�:���p��>E�JuY�p�*Cʇ��;�`JLz�4�e:2������˗Fb<�f��+��J�W�UG%'����j�����Âq�l�_�τt��@ς4�A�5��|߄�v����61��Ϲ+7�[�,���Ώ.�����}5XA�)�X���ޖ��4TMWу��d�2?3.� j�!�9���~+n���rM�MG�#Z$/�¢	cd��6�}�d	��ȟSd:1��l3fN� �d*O�B�f�sC��g��<�}�=�����^��Ct���]�'��$d'�IcZ�3�ӧ鑓��nر��؊@*��i�5YyrJ.]�2$��1?��WJ6��C�xoz�qxO��-^�˭^>���U��d2�!��ݿ��5�i�իF�'��:�fBWE�撈����s#6s��:!�Xh���R�!4o����I�g��5���޾oW��"�����(>��F��=,O&��
�ݱ9��4(�t6���8��kO��}��l�뚖���B�T�@�I�|�>}d*�HUd9*�9�p�ԂE����7�^>�z�u��m7�7��;8��ksD��%����B�Cy�90�0ϲd<ռ�X��A�3�v>{��1�aEw$=�%&�S�o�:mW�b�:zs�LNc��j+����c��e��O@H�Xi�8��c� �W�$g�9�#����1÷o��&r�A�.��j��=g��MV�tSjy����ѼC�F�/�b�Q�W�@��Gy�"�Vrzώ��Y���*�6]#V�a�G���nP�^熯fl�(ǻ %��!`K�����"�{jd�Zw�8��xr�����
,����?�ԓho�F�rwc�4�c��Lb+��F�P0�[��2�P������M�����>z��|�N)OJ�eM����7�E!v�6�S�̕�#�;�/�q��쌺��}��Y�v,p�W�d�R��F��x�_�V8+Qm�WD��>X�*�wI��R��\ϭ�}𺎌c�Mu��2��c���n�L�;�������HQ�Ik�mS������ғ��*O������:���d�oE� �OǷ��'?�gd2��[�^���3�*i��lk�G���F�҃S�\�G�L��&�ۻ��u) v��h��f��+�T�����o�"F�_�ʤO�	AP�v����<�9:�wk���K�=�X���@�ުN��{��`X+JP5���ϳ���F�9?�U��a�4�R��m���f2P��Aek�0]�"z?�8��044����t��s���93�}��'bz��!NB��[e�zN���X��7"߂NaY�I*�Vj�c��i38������0�ct*���4��s�J��a�ݮsq��'��}�3���vO����C�BJH�LIP1�*OO��ARt�oc�յg&��X�EO��}����%C��dD�Xi�ዪI�|�lK�ڷg�sĺW�1���S,�xk ,X���,c�ޥŦ�c��K��=����a�}���4Y�v���T��2>��7�KX�iD�
NV��ED��02S#u=�*���Ao5���� :9�/t�����u������}K/��5��y���U�L�mt�>�K�5��'ℸ�N4'3uYc�d�г��H�rAv����9G�0�
y6�he���:��l�Z���?l�\��1�R�a'õ�(�������-WD8��̅�8p�s����dQ��-���G(����5o�����Qf��]n�"��p�7q��:g�H���?YK4i���]�4dQ�ץ��U1<��;�G@�d�x�_�6_M���'�V���r�e�����_���#_,�i���5�N��YGWR��?�O�ׁIVeW�9F�s�<mo�#\���&e��p�W�^���ź8�5��כ���CR+$���k��y��nWx�p��S�i�����7n���A�g�X�{���g��5j�����C��	")x���H$���[+%됐M����i]�%�q�j�>iꭠsނ�<��HV��OY�f�#$d,H�} On���Y��� ;g����U�ae�,�A�"�I��՝���"��ꉋD^�6�;�_zeF*��r� ���P�9�{��� L�F�$�h	�G�N/VH������%��I�^A� ь3>%9���^�;��&D(O^Ȓ�����x�,%iis�������?�elb�5Z`�]]u�[�k�N4�YwR�I�k6�Yp�C�%����$"i�u�����G��?��ҷ[lւW|���. ����Y)G�6�w�/��>�b��5�1�k��IY�#�svA3��~3��5�'�3@�_�e��!�G����iI/�d�O�
�w���j5�	�~�����'B��:�g�gB�;�u+��+Wʽ����T��%����ol�q{!~n�E=Jv���(��۽tٗk�:Bo�^�~o�*"�mL�W ���l������z�0_��ܻC�̛!z�sn��iV�C$3�Q��!f�+ -�ˁ[�d�Y���|�FS����7�����Ր�>��vv[(�l��A)ØL*�]�������&��xRnC�"]N8�N#F/�;���d�,x�B��M��Mi����M5w���(�p����ղnR�뒧U�+yD���::|,Zv.�h�ic6ȱ��v/�(��z]7�����F�F�}N�U����A=ą�Xaӝ�J6������=d\�����-��W���x�]�A.�-�1��p��Fr��-n�0Hb�Ͻ���e=��XԀ�|+&+ł{84�<�6�Q>�#`�m�3g��l���G!�Q�U?�e]o��{���@��a�+�e�p�)	�L��ҋb�1c���0�<�'���=�I��뾥����;����^��U�ǖ@��U��О�,'q���k��t�J� � 6���r�v��6 �O�&�+lm� �lTvqb.�s���|�<�����"+�Y'���>�W\�o@��0Cu�[�d1����<������q0b�����-��?��Ϗ�E���
�W_���ui��(܅��"��]�n��
��Ћ(&�/5U}� ���?��Z�?��̙.jP7J�}3�x�ţ�طKlA��m6�9ѼK��d+��6l:k/��hE67ѝ�����QY+��6ő�_��MK��_e�_��Q���j,����+i��<"@>���P��R�t?<wφ��L|UkV�	Q�Fу$^# w沼]���CJ]�Qy�U�U�	�Tͱ�>f�=���J_���~�e�m����Q(��Л��å*#d�)�e��8q�7��[lϕV����b\���%�s �"���/�:L���B�ܣǏߓ��:xj��>��_�?���Ri2�W�&�|�֖<\H)0FGy*#p;�xq��TE?fj��$"�����#
L��|�et��4�
E�zص�f���;k�ʦ��yy@�a�����"��X��y6���	�,:9������̼��h^|83C*���'
Qc�˝ԃ<�S��W�Tp�d89JL���#sޯ�C��Y�G�_���C�Å{'���!g���Wa>PӒ[!7�Τk[�s��	Ǆ31ѣ�%� r�4"֖�%P}3�4wo�@!OzSn�t�?jۦ"��!`�U;�Hٺ,�r3'���y��6���k*�Ȑ����� �N�����o��*?��V�K����&���"2�>=2������x�ꂝ�:�'����T:Q���{�i�s���;!*�ź���2;;a�E�>8���tV(y���S�#�v�N-�Z�:�7O� ���E��I,�ԆUN>5��n�U�١��F�w�����s��Q�����'|�r��l 9\�=�]y�5�c=�YsK$�N��0��݋���ħkn���B"y�77W��ߘF��2
�,i�5ֆ�*���Z�*�<߄��0}�Rcc<=S��M_�c�y��U$�e��v�}�����4,�ϻ�ɒ�pB��c�u��+ƶcw�̀]oKQ��ȱOUQ��d�Б�/�5O�N��O�.V��ѯ���簯28�Ra�Lb��ֽ���W�d�*#2��+{�+h��u��g�!y#��;����h�#�Q̖4<׌
F.z-we�>�]D�)j[,2a�0S,�����"�8��������)t�;����8�	�J�ؤ'�{���84��{��4�X�:u}����@�7�`U�2[�7F/��/��,|�M缀�F"uK���x�Q���� @0�Ǭ���2K9��Tj*���V�{R�!�X���Y��{Fr�}������҂9��z����*m��'V�u&O���07C��`n3|Q�JOQI��L%�᧥t�~�H*`��Ah��~'�߃`0���Eu�Ƨ1��v��B�y�l� ���v������Ij��&���:��V �AV�D�P�Kb�2��z�"9$�����#�l����T����EZt��n�:�O�0h�W���\}!�W��*�mXA��@r�0������߻���,B߳��G��P��\�U��_���ܝQ�p���Q(�LuF�1];��'��WEK��M�u��� �o�Zՠ`��=tt�&-�o��w�k�b>��ԜPQ"�V��N����gY{��֧ؔ
ȧ�ﭜ��%�y�5�LNe޻Lbx�M����V��qs�������Ѯ�۫,�Xюcok�$/�����'s��3T�R��Nx��Z��<2w��һe4��G�᨜����JWE�z&o���ס������<u�-g~�S�w�D	�����'	(�Mb�2np8�x�v��@|fO��NM8�'�9�Ei����u�f�\u.���u����M�c0L��3���\�\��aw*��~&5�`��`&�X}Q�@��)�ܰ=�J�m�b/�-?�f$Ɇ�є�SYVg��5�V�Ƨ����	�����T��W���ط��9�^K��\����7q�L��TqWS�0�9��]��6��~f���/���t�"":��.I"�dl�[�J$��pd����q�b;��[O���&Z<׭���&���\�L<�\�>@ՓG��O�mﮬ,��7���Ń�r��L�mFb�X��n�+�L}:�e5��7]�]k��u��;��������78��M��A��(�~0������M\��׎WaZ��?�k�C����%�S�������j�\� �e.�A�ͷ�KN�^_�?�0�l,ۊ���?4l��;��s�������c�!ǖ>������W���46�d%%���6F�M�?�=�&��GJ��{�%���m� oY�+u��%�2���ލB���O��1/�,B~�8>V�ܡ�kVZ����y�I�jnk����!�Wu���Ti�l��nz��Z��UUAe|���T�iw1�����ޞ�&��G���@�W0OltUb^Pc�0�;̺���:#kC���ix�f@��&�um��1H��������$� `�&'CrP����	����4QPn��14;�1�<��w�;'�e�=�`��y-�����-�o7#� �\�r�i��b�� I��b����eD�W5��;9�s�����EF�GM�� ����#� �苩F���w�\%�����.�5	y-����l��i�B�(�YQ�� ;�c�����l�bu�ȿݾ��Ǯ���t׼W�s[o�m�J
���G�6��Z*���EZ�BάS�%%	N("�}gN���iCEW����J�O�c6��iK ��E-�����|�P?�H�%�$_ѺoH�w!w_�R5�!s�'��M�:�&��`�D���VG8�$��{ �'����B���W�.m��x��&�T�3�I��)�ÊHg�;>X��/�M�
��7���Wj�[����AE���`}�${���DG �����]��j,E"�����}:�R��ԡM8��w;X#������]�g�Jb%�:dٺ	E��� �V�e-������M����z�����WM"zl0�$����V(�~��!S-f"e]�q��Asl �}R'łO08ZJ1ʣ
���^�h�����!�*���#�s�-��R�o�껡O��1��BS`��i�Z7\W�,�h�(z;Y�/(B�V����D����~��O��^�C����Jt��H��`��^�UZ�����A�vrHE��:��*�Zl��=F��] ��r97
�{(��80�U����׬���2+UQ�,(�dGlpn��Q�^k��V����7�)���B��Ƭ}��0�I��L_qBṄӃ0�!]���Q��<��)c4J�\D�ښY��
�]��{��&P~vR?�u�hf�/gw�>��6��e��i,y����O$�����?�6��Hx���7�۵�ՇYf�(;�Ʊkrb	��3І=��Ё���
�1�f�s�N�+y9nͬ=��jTTEh9gNs�:��Y�>��n /�rQ�`��ͺ�86Q�m�O��F(��,�abS֑��W����Z�2;�@�M��B�oL��WP�s���HkH��Ԙ/��]�;�)F��DA��w���ς4�R����>J���8I%vU�\��tY^���������T6=:@�貊<��ޤoD
�Q梲����=��\������Xw�n��yb��{��[S��X	��<Z.�-Uk
��h!�4Zχ3y�Fo��q�㎠G�[3�#���+m����r��g���5)��eu[���׍�O�{��˄��ǭk�H$N����=�h���SA�p���x,,���'�;�S��o�mIɕ8� ����^��I"*�
~�#��`�7�K(���Y�*AD���sީ:����B�Z0�K����~w�~w�� Ф2��{g;N���i>�g`Mm��d�~�������W�޹K��2n�Qb3<����687��v!�Ȋ�nǤ��(����@�W`ʸ6���ŕjl3��U�����W���q�*(+z�C���^�I)1��iQ�,��9S�����7����?�6�iJ�L&���l.���J ��IjB]��Õ��,�0q�4�ĭ�3�.-��������ae
DX���$�-ޔ����^��&���Bsu?�Wʦ˂�a�ll��Z��vL�i����}��J|,���?,;UA��DW���^%E/���/ l [Z(��h~d�=7��1�zN;%���u^KR����>�;d&�S�UVi-���xlJBW��S.�1��NUR�s��9�'Z�C�F���$��O��M�$��V!�jeEH��9��VHܲ�%E���[2�nR�ʈ�w��	@4b�����a�>�n�hY1�$y[�>�����V��$�!�$QBv�2�2A�rkT	�!	��Zx�v��W��W�f٤{O��l�,��������M{�X��z��T=������f,�}��Vc�/]Tb���	"��O6.���nv�4v�93��m�H����O;�7(MBR�u��?2҆+�w9��`���x��T����z���n�bk��m���}����v��`�}km�+�HP��ڵ��mbW,�ųQK����VΤdطC�~�1�й�z�u��2��#u|p��c�E
�L�9@磝_m��!2씵�s�7ǒŋWA���n�qw#��,x?����t�N�}�TF�pi������A��U��ʳ�74s��g��o�	R�D��R��]+
�3�}v�vG�.�KRTl���D�:77{��)�w�<~��j]Z.Ҋݚ0�t���^�^�"zd����	�������k��F0UdY1Ɇ~�>���p�|�b���R�goRv�R��R�h^$˗2��6�ȳ��RQ�س2�L�0�_��l�*��|tW��E#�S�ÞX�:����#�!ǆF��Vwl��&��[��uqd�x��kU�Rk�m��1�W`�ˊ��eww�E${`&隧/��	+zm��${Qa��A��qTζ�߿��Д9��*9����'gH�_��@���>����"Tb��E �U��܇�J������#M���D�3f�3$�y):�O�qh"F�lo�5�(�� �{wD�PK;q��7fN�@{���h��첏ަx�TO�&�So�;��_�����[�L&aP_ҰP$���{��p�E�fr<Eg�x�VT���]l��D�����V�z4;��pi�bѲO������dβ^�w��{�hrm�(e˧^�ٻ�r���B�7S�~Is�I�fό����{oH�ʵ0[���?4(y Z�b~��m].ت*�"|�����C74]��Sf�ZB��Ѡ��j���w�7Hϑ�`	���=�7���e�
*-�H�l�l�P��}|��|��ݽ�c4w���]�e�e��3V	�S�d��������������U�gz�w�o����S�ߕ�C"��?m_~�F(3FlF�9��{��Bf#��� 7�_D]]�km�/N� ��G�����5Kn$�M??X��,m�h���ǆ�#LQ�T"��$2u%��W��E�¼3;��%���O�>�}�]��Q��k��rU�w�~�ݿԠ#�Cm�&�΀�gb�B�N�ޤ;�����
����+9��)�T]:��pt?	E�q؈?]l؋?�!��y�/ߛ0TT�c/���^9
�����R�5�n�ry1Mcǩr�z~,>��u�(7@���.���>>�.�>dﻁ�s�A��ό������;GN7�I���x���(����f�0|�Z����6��tP�d+�9��޼��`1"���_t�[���	N��-�a�ￗ�?*��i!At7< �_���C��"#����6�(��Ձa�o��,K�#�b�_� �s�P���&^ V���� J�R�8�?.��n_�D�
D���h[����{�W���[���h�J�*��Կ��9x��P>��-\��rMΨg�,�~�g�$^YG�@���4d�(�g:�@��O2���8S� ߳���ë��9]�L�=��C�Ps�>%#���w�h�VV�$��p���ҏ���ύ�����[:E�g�A��qf�f���}���ݧB��� b�@t��;2�b����m�'���e��Vf����C/e�S<���B�p��`����'�ϋT]����i�y���+J��X=�:1�������6LG�?+��ڗ7���p�QL=�|�-�6~�Sa�}����?h��qh,[���T�S�QW���Pg��|~�'�ʣ�J�������q�M�I�c����L/�]y��������ǣ�K�ZxIk���'/�����'�g������ߔX_��&Z�Mkwu�i9�;s�JMG�K��3�{}&�EcZ�˃��	󗲏��v=Z?X3���x�7�o	B~����d����fvK�o�*���n[��R����29�4����df6�hl���r�14����	����'�(�L�sm��:�&�l��it������k����v�W.�|�,1:@�y󻚊�[hY/ð:}�k�m�ua�r�ע�\Ӽ�O,]xb>KM�͸ߘ>�qg��4��aW�;S��nq����ܾ��6��D�H�Tu��F�*�_��sA|��N�o�.��.�!!��;��LrI��� ���q�B��ɺ ���<u�D��<ǘ����"_
~`�>�'"H˭c�e�$G�W�0)�Ȭ�������<Öz�u�����Cu3мΰ1�Ÿn��5���笍���Ź�h���w�\s<�v��C���_(�]1!3�U����nv���=~�����b,EU�
�cDg�
cIP��"���<�Z�Yu����½JN*7���|�$�Pr��1N�����\, ���^������4X�ZO[k\7~����cT��|��{n"4�v�I�'�'�����ĉpn0e��y���XP����x>��Q���qi�/Ђ����d�Uv��k!�_I�kj�?���)xH7_¹S\ëU��`��\�p����#/�Eg��n1X��3�e�ck��ԉ��f�gic6��.ٟ2݉�����]����7�(k+���S�l�fΐ��f���s�N����	gh.�c��޸h/�B��v�s��WBw|ǾU���Sx�h,%j�^��~g��Ժ�`ڃaRlͅ2��;D}p��������ɡ���>��.�,F�v�)�K�i�b�%|��Q�2e�f��	�z���1�������r�DO�@��.Ɲ�Q�/����⿭	��}x��nni���lY�*N�	����]4�pt.e��3�/!���(V/��n:�R��X����1�K�����#����B,G��d�`MP����4CO�E��C�
����J�6D��&�{7�������pc���4v�(%���+�Ldx
��^	f��,V&�^�{ɸ����ע+'8.�f�ܤ;K �~�Wf�}�W�g/4�;KQ���[�RH� o����<�>��c��H���u����o�d߳C������N]A�P3#�D���'�A찌�������W����]����Pa=_hh4nf���I�`�Zh�ë�+������nC�>+�н�?U��C���N"c��JpZ�5u0�Ĉ�(�1���+�*Wxx�g�׽�A�Y�Ln���K��K�N�i����`��^rd,V��[%��ĕ	�串>��p���)8>5��~-��`�[��_(R!�!Y�G�j��.�
�������&lдzq�P�������H&�zЕ�l*��o�V���B�W��@����W? i�D�ME�A���*���9����T��U���u�ش<�B�	��'��hT���tV��%m�0w� U�� n�	�²��:lΰ6��}�>��Jc��P-�趁ƓPQ��j��24;<�쿁����Y�uN� �6�n2L|��c�Ze�������OyJ�I���u"�c�N�aϸ��W���
�,�(�Qe��9�_=�7�����X�	9��������r��w��o���R����)�ܥ@x�z���J̐uxn���>�&�«��_���Q���)�T_'�����,d��sDK>����zv�ܛ�n��s�!ӱ���V�Pgr�����b���\1u���*������E)�A������ȹ�öZ�v�
�wc~�����x�jpY����G��]Y��5ٓ���=�dӒ��#A�_�gWʻ����p�\�=�~��[�B��xZ_#��\;�局T� 𭀓�mr����;��"w3Ȇ�&����G�{�Κ��vS6�=��!�D4�uY��8ס�/8
�Bk�ˀ�"i�C�e}��M1z73A|Mf��ҰY�z�@y��nc��~�¶� �ڟe�o��<s�|Cs*����r���"�۷^tS����3����&
��P�p��DHA�yj�'��W�َ�/��
R#S�F�t��b�MP�L�Ȭ����?�ݑM�%�>��B�-�����~�:��Y��CFݺ�'�FH��m/���&]�cK w�4L�������c ��:��� ����ox��� �c�l!#�}��χ{�<5YPk���
�&tU�������.*�O��*���0�����G2M��IPd���H��@g
�BJ�'V������d.��o$��=�V�H�{��9��--~���5��p�s<��OA��	�%=7�T����T�Q�v}v̄`"����i����.z�����UiJ�w��(«���q��� �a��]�*#+�Q-��Q���uZ��� m{�ؐ߉qة�i�������:(�*x�j�b�|&��;�_b �����豙9�R�����qx�a;a�추}����s=�{����x���4>��&�G�I����(t���v��$���?�J<A{춤�7��7��YH{��.HQ��y���O��_��قt�������6��%D���1��'E�	���]�
S���܃߹��?�Ci>4W�Cw���rg^��xڣ�v3P�*��LD3����������{>S�Z�ڙnX]��xb��s��Q�V�R	���a)�-�[y\����B��뒔�^��i�ِ=H��PX�
֣���/�|y�L0��#�h�ɁkWf��<�Fח(��SRj%�|�yø6��w���hc��=7����Z�Z��/���.|����Ԃp�-mݝ���:0=I (��D���5�Ѝ���#�Z&~x��_��)��`p`��&(Niݧ����w4��ܲ�o=��9�����TBͧ��o��_�� �Ss>�Z)&�+�Q��f@��VN|��i�a�D���w�A�~*�-%���f�q��] �㷂�uSw��2�ED�+���Rv4#���y�VD����s �`wu��Ai��ϱ�x�8^Tkx�B��&�=rө6Y�hH�P�F�YG�U�$�Z)����ۍ�.��gO����.��ʼϠ�5�7�͖2R�����k����n����?���T��=��h[]@�ր<68<5�y0���H}�a�ƿ6ȱf�����z���_����y�\c� ��:(�2r���/$�Vx0#���Y��ꚴȹ��� �:��q��\%,�|*%��.�_�S"5�����1�K�f����� ab�z�U�w|*�� �G8�u>+�?G�]�Х6H�)��/$H��hOp��tZT��Xj��Q�OQ�rȭ����z�~ss�|E&YF�m��}�R@)�3`�+��F��C���@�A���x�J������o��؉q��5��U�.A�,���O�8�����kL����u��tR�f�C�9�K����Y5Q��f��L�kf��%��,HF���'j?��(�+����JI{�����A^̪�:����>��'�E���Բ�SÉK�s������0���H�6ۏ7�/����=�~W*{�>�B�;z*�?5��zq�v���$UR����BZ�d*�S�(�E;���=�OL�`^�ߧ'%��A|[�V��‶��O�/��������>>h|�s�]3w�i�o�\9:m�&y*g�TПL��ܠа�4�M�v��&��lt�;��XP��f�a�j������t���X�r|$_�XR�3��y�A	~�k��I�˚��g�g0}���ᆪ>�ϝf��#��h���1�4�[9��.�,���c.q=�cQiD�"�:pݹ�Sr��u�6�3���n pD��DE��8)6rt����'�p5N���ظWt��ҹw�?A�6��ā=-�#��V[�>1Y��q�󠎼�Â����B�u����v�-�3��
I�r�Ӯ��[��*��F��#���@�~�x�P��R�/T�d�����10�=?�� �R�ٓ����I96.-271qH�.�vJ`·v&?��{�s2�����ʘ;XW��JR
���L�Qv1�>~8�B��\�9Z�38�Q 662��6����(.�c�\�|wV��y-��1n��8���G�e*��}b E�u}�������eϞ(�L�Cς�&�!��V�Д�tg�n���lĳ���,�EJ�YJ��v��J.���v�ƒzD�����P�q��<�w�|I$28gBf�o m�[���פ]f�P��l��ar�n�ׯ��-���ySnG������M�y5Z�xGZ]-�dP
<s��a��B������tZ�ݙ�w��x;�G��T;�R�`�dW�˧�ܮU�O�8T��i6���ߕ�)R���E��(ʺ�&�>����o�
��A̭�X%� �uϩ�<�)�Y���a��U��L
��a�:l7Q��Ɂ�y0���T�n�0E�����\����t#������k܏7��k'��K�j.ж����?�Q��E,�B}H����&���� 7!�C���ă���]��Etg���7;�)d�ڠ�"�K~I����E	���.C�l��,��@���;�����&����K�8�]Μ39�� ���~T��?��mOj*��hYMڴ��Z����(5���ff�i���7�߱���F���e�ܷ�;>1�����\5c+�_���l��eh�4-^�O�#��R;��MM��,��8_�HߺN���!`���8j��T��N�$��� ���WAk�Y�5�H4�M�u��Ű���������Kdlԁ��R���|-i��p	����4�x�q���O+��s��Ccq�،z8��T��h��3FpP��l-Rk`bbҎ_�VϢ9���~�ف*j�h]@��i�M�����j}3i��.�L�⍸ۆʒ��g���?R����
5�F��SŴS��G��&s�%�؍��[=jHڅׂ�f�%��`��:�V�(V�"8T�s�MA#l"�X谵f�hE�W�q��*`P3Y�:vtkr����x���RvxL��������Me[�����+�s�+2
�� ""J1b(�0#�:��A��Z0�6�U�Q�9�HW1 "E�^"�`��[B@HI�PB�w�s�}�?��|���|��>k���w���0�E ��b�>���f�}�J׌Ω혢H�����"�(�=;)�B�OG��h���[�ƾLÕ�[�i�e�6��!Ơ��LX'R�����L��*���#[ ���(i�@�M�Ǔ�lI����w����*It�2���_,�_qi�������w��_˪�峁˼(�+G|4G���>�5ޠ�Z�k�뎩��ʾA�6�IO��K� ���i�چh�S#1IJG��$�3����x��;�3�f�~�;�H��o�鿁3Lr����a;'�Ľ��X/tLU�:����N���+��A<����N��j�Hc"?jo��\[d	��mp��F12<0�67q"�b�%�)y���|�&���
l�ܨ=�լAY�B��M���M�Lg�OR�tZBC�5�W_��~B<�;�ݝ���oz�����z����K��i�m`��k��ȇhّ����� �a^h§��U��g��g{����7��������vz�ޚ'|��� a"�g���`����SV�L4�Z�b;��]�m�c	(T��г��l&L͛Z��V��݃ڪ��Y���zk}��+-��L�Qj�`��Us�����=4i*�ܴk�L�U�;��HC�Q�x�4Ӹ�O�<��w��ʑ%hr���HΛM̮�>% �䛚����Ԫ��	k�k#�3Ea���O��{q�~;�Q�0�-�J/V#{u�����K�}:�+�%vh���L_e����f���;n�(�3�f�F��W�����������Zx�BWؕ���f�of�q���Ӓ�I�v/n��[%՜/�ܨU4x���R���2�gO�.�G�R�p�ގ�q��)�6 �kY����$٣��#�/b˴_�k���c�������_����HTF��F�<cN�i	��e��� &r1�Cqdۼ�5n���J���7��ՠv�k]+4�_�q�ablxX"��Z�Y�m��uL�&1y��^�r<��Uk<NtZX@��e7������ͨ`�V'����˦ui'�xy}c�s.D�#.�@��U/�g��h�$c+ҋH wt;�2�n��U6� ����|���z���楳"i���3_U�a��ZV��\�Ò��K� ����v7jxdg����L��5�@�F��U�p/Y����ƍ�S�x�4���y�7�1�}�;�7�c�t��o�ε&Id��vSb����;�ƀy����x����ܐ��dgb�a����2Ȋ�[3%��W�v*�x��-�(����o'oC�ܷf��M��N���!�ԥ�YX��")��f�w�:�e���r�pc5�#�a��������u��8R^0lQ��ޮ����>8)H5T)G7m�
5�o����3y�aQk3c���#��&�gw5*�3a��S�޾���Uʈ�a��S6;�[��ns�@U�Bgc�����EbXf�� ���jO��[|%ju{Be�W >P��p�V�G�[;/s����*)]o�>������aL[y�
����{���4�s$AK����c���g*���Ab����TI3�$���$v���.���x�Ǉq����j�"�X�&;�Z���1��=�`7}k���p�P%�=<�ȕ�{�Rn4��|L�$���gMX���h�`(P?����-���G2�{iG��R�?���/��쎥���4�z�_��~(a�%%xCh�`MIG�,�7���B��.�"^s��h�w/�[��4�e�~s�Ɩ"�>�5p���7����kヮ];A�IF��!�`��3�񺒭dT�F'Y�2>����SV��Ǐ�ێ�t+�R#�k˛ƍI�����7�xc5*(���|����ONĊ2%��%��ȿ���K�c���e�SY���rT���\�U������V����"�[_�FӱZKY�g:qhs�+P8�G�
����Qb0�5dP���2�C��Q�z����&���|�ٶ�~s��iw-Xd.���Cp�B��k�y��Wg�z����A����T��3��+F0<��E���3�=�=�"U���� �(6����d��g�>5E���t\� m���;2v���"@* ���I�1��4�	��U�?�Y�˨�G�����*@���a��%*�O!��v�U(`I� і7kh���v�T:�ٖ�g�u|k���l�\,�3c&��x[Hh+_Ur��|������������H�L?#�3�5����mc=
�o�!{���Y3�/*�GN�l���	.��=|aKC�5O�kd#]~��6h������NjD ,-F[}ܪ=*�V�I�A�Y~�]�ۡ��6Ho�@)ϊJ�e#ms����w��є�̖�ϽiM~u_�7�Q�f�C�s
Bd�G�J��̳�1 g�q�wO��湠���_}��6�\�ffY����ؾ��h�/�Xgě����E��,]ZPp�-�@�� BmF>�%c$�j����ѵ_h��dC( �}���v�(g<]��K@<HZC�]뫵uTmP��NI0#V��D�5����7�ۊLTȝ[$��ɜǀ��
iO��%�^� ��oղ�0������.��h�%�'�g�Ɗ� i���~�Y�!�k���7;��� 
 ����Av�c��
�8���N��ϺcE:���ϻ���1ό[I�K���:#i,����My��p�v���2T�Yß��o)1	A��aF�������x<�q��(kU�7D�V	� �M��:��D�^w#�0(r���O�,���j@�
��0+�����
 |��i���p��f�-�E��J��Mɍ��K0j���C��~f<csb~,��xDŤw��1%gp����gd��c���y��]P�2tg|��b���ț�� Y�S��8�<i��M�(��]��x���.� �ŌO\�w:��AO�� �?���h�2�c��w�wu�H�W��3�Tέ��{�] n���rݿ�a	�O��*�~i����|9�>B�#�La�z>>Hr�!�q�oܛj	4|�|����sv�d���#�������J�@́�����;ekm��2@Bu<FK��.إs!��E3����@~3v�~��A%�0@�G��#n�(4�k1H�*�W�Q'@G�yP,&�ghj��3 �W'y,���2����Qa�MĻ^�ѕ�d�F�����2��a0H���#�Z���}w��Q�ڋ�i���e��n����p��砀R[twl�O�xf�մ151������/����e���6��d��,��T�>,Z����{A�}�?o7L4�S����� ��u���Vgu�����z)񹒳#�
��$��Ǩ�mFM��ۨT3��1��o���r*B`�ǩ��l�9� ��!O����b[=�\;�(&v2݉^)�-</�"�e1�E\(��}����S�&O���E��)�\��m�B�  ac�u�bC����7`��Lb�)\�=#ǣ��81\W������� 3:f�Z^9�cw�[���� ������6,'8��+-��r��
��pQ>**�����
7��,�+�kw�w*/��G�K�` ��"O�Z�zP�$	cq��V���x��d`
�]����]Rfa��LE!Pt=x����Z�/��s��-CI�
n$$�B�� �h,ù>n�u���z�ºJ���	 �v"�!�~6LU��^�͊�%��Z��K_ *T=��b$/x0�0�?�>Kќ����B �M'�T`H����j�SnL��8Hl3_�>�m��7��t
;�a�AdK��}��&�z���C����r��n�Ҝ��{q$��9� �+���\|�
c��ٗ���`�^mG���<ި��"z���Y����N�%�\����>���o�!��?�pZ7�`�ô��wJjn���ܻ�9�UL�X�R��YR�_��:���Pٖ|y ��t}�i������F�xC�����q�'�C�Ca���5|�O��Z ;K<Q9^(1�����T��W��y� +3�e���t���!�1n<�W��Lu��v�!zwl˨���2�����Wq�z��F���3ޙ�� �s�,$f���+ ��(��oj����y�W�	�.��Y���#xw�Q����1�  O�C�;u��tl�(�󭻘�9�co��e�j�T��y��1�	zH5#,��ɡ0�IF|�s�͖�ɗQ^�����r���n��@����o0�j/Rf���;Zb��l�c�|vm�tc`�P\/Ā��]� ��!Ts�\�'A1�� �(�x�S�� n�ѓ�1�?�5�0z/叝�����|���a�X���d����L��f|c�z���8}��������3�ȗ0xL3^�"�m�$�c9F�=�<2
^��5D�eay�I١-�t|M���v���q�Co�z���շ_}�������_��_����o�Ҿ��+G������F���]Z�>5䁕�����__���չ&iԯ}`=O0
��J�7�w>v��|U~�0��P%�g{F�Os�xGK�D������ݮIQst�=�]lί,?�28�e�ш�F�O�v_,<�-N:�̰"5���[��^m����C��aO�۶�a���N���A�5T9rW�-϶���}�6z�®X\ά_�x�Q@uqĽ;����9����E~�3v�J�OB&�� BnYYF�h�R��r�|z	�E@��_g�i��-#?R~p�O��M��o���Z�0��@�ь� F]�	�����6��%$����~0��O��Ԩg��*��{)�1��3UF-u���»:��L��	j�iIl���~�HI�����v��K��� � <����u�L{8��W0��q>�	��a��!�'�D�#҂*��@�,O�v���9��z ?F���e�'V�
��p]֯�?G��,�\���������ǹ�'0��a�q��6�������x%0o)ݺ4��S��t�M2o)���=T�O��G�+��zĸ'˳ꍨ!!e�0�cN���Ӿ���*�J���)#�-bu�ܢ԰���O�\���T8�ed����h'c��i�>��v&��;�T�j�+�k^�����[C?�%F�/eK� C�tU�w�BdBY~����+���4�YC25~^s1�
_�T��i��1ة �efh�?9OO��z�u�%��|�?��nO8��"�ax��.U1��y#YG�ͱ�������R��XF�G/T��H�ϕ��~;�~�$�1�iL�Yܕ�u�X@�g���ZUG��eU'M��? go�o?8��t+v��E�@b���(j��ä�'�.�<Nh����3��gB]���	=�>���}���U�Y�U2������|�)����^4���{��Vo����VVgq�FvD�t��O�:�T`*�&X�G��ʱr��0��LO;U�>I k�Xl��ʕ� ���]pWb���$�ID���Iv�i�h7�C7�U�"�p6�q�w�U�S��Y��F7~�"g���4�rgUݵ1��%j����C��1�y�����9������39��@z�b���|4�Ǘ>��er�G7~��� -���<��q�9|P�kݎ��Oһ�:�{�ʮ���#���B�V��3��/SaǈbdiA�)1z�B�&ܔ��V�6�{��o�d'*���F�&�7b:0�ڦ���akW����F*<�ꋿp�j����6l��ZL����(_�3$�ߩpZ��q,?hߓ��KH^o4\��IY�n�$Ͽ�ɃG�0r ��8+ݎ��uv�?�+��o�h�\�R �_K#�N�-7���"�^��k��L鉹����e��>VР�0g���Y~�)7ZJ`�
��<K�|(����Ȗ��퓻�\�b��d$��ػ��s�m������1h� �T3�F��y��k2�,m䫹ſ8c��r�ȷ���i\��j7 Օ$���n��B�D�[0�s'oIVC�IDH���
���7n�į�ni���շА�K\Bn�E���Z���b"�8����[���[�A�/	�V��;`�U�������ḱt����'Y�b�\w�f(����1m�i&��ލ�(����!�dH몥�[~��	��[C0�*Վ��A��pȚ{7j�<x:��(HHu4'�[fP�~Lz���P0v@;"�2��G�4ǽ��цG-�~�j��F�z���.�ye%�]%�_D-�F�7_�ʸE��d̶j6]�@2*�O{lh��y�\�N�ҝ��R7Z��ep���xu��(�t��e54���@�UK�2A��1����]�	�y���o�^�*��D����9	F�Wj�Ѩ����W���Q�D��T�	��	��8)W� ���;�6�6�
0r��lK��s l�ү���`�x�Mo+��,;��,�ӊ���w��)��]��F|��]�g9�C�+k�J�8�B�jA�Va(c�^`t��>9�5'
(9_}R�|2z�tX�o�Nk�- ����ֽ��{ҧl �`u����ͬۡ.G�^�eȻ�6W����O���7Q .qK��Qi���e���b1�Ϊ�㣖A���������k��I�G��R�I��f�>�l䀉/b[�cG���b�C��O�����}c�]��B�����1y�BW��4��a��~�6';���տ�V%��EMk������pR מ��4�F}�q�v��������/]m|9��55��YD2͎��$IF��������2�Y�VB������n+�%�ro4̑2����)}u%B�"�`���a�P�����mkX�Aއ2�:o}�������@������6e�ŧ�ڻjX��Q��v��ZH�l鮗|'�Y���)79��5|�~RN�%�7����e��Q4���eTȁ�n��F)9��h���!{��^�i>��FE��&w���G���mW�u����R���қ�U�6�v̐�����7Fv cO��M�H&��+c�fA�#���~�J��T���P��ڌ��Q�<�i��1�L
?�u��A�(%��^_����$�q�z���[��&�c�`"�e{�=dp�a
"WZ���z �[H�ߞ=�O��ظN�\v?>��d��<�٩ۏ���#��N�;� �P�:�H!D{�$�Y�HT8JO���	�8�j04�Le^��E�J�<X�c�R�$���޳y5� e�sh�����you;�|��'nr+����;���q�9䭪�<��1��Z�9��a� ��>i��#\�˔��`DR3��&977j@tҫ�k#�*��fk�ֳ�s�_�Go|٫$-h\LwT�	p�yX�{By���v�M��BVw�.�k�� �������_��y=4������u���%������ߊ@�H<^5(�o�2�0��՞�)�ҋa]Y�j�u �&َ����$$�4�Ƨ��[�0	��_&��`hq�xr�M#�z���uO�(��2>=W���U��J����^�<�>B�N`�aV�����W}ѻ]n$4�GG�|.l|��8�s?f���럚eT���SO(US�,Oc����2�FƁ��@��0(��d�ضn���v���u+��B;Y�XQ��	���_��!�!������g� �)����7��<�W���P�h��(�4�<ډ��hz�F7���=�D��eKRӄ�.^&�C��򋻋N��`��矚Qg��*'���׌�1�%��*-�Z�ږ��J��'9���-�1���v���:P֨�:XY�=@CXS�xC4��d�}���1� Ð�����+ulA�Y��J��hEQ2AZYv���l�Id�䞨jF�+ǻ�!#�~)� �ƛ�<M��zK"#�X�2ΠM�t���@�ȣ�Bj*3 ͜�(��p��a�2B_�R\]j�;p&����䟠8r��1MU�?�p��m�dB��)�G0�rn��ܖ��C���C���č�v>9;���v���(�~����٪V9*vE'�D�Q��z ׁ@/4x�B�[���ض��q�@h A����{�Te'Nv�Y5�jΧw�T�A$�q��0��(ޮ�%�3�����+'���b�;n~=�q��$�Ӓ�o�v�[X;rs����E,�Ez,Y��5n����_�|�9J�܄�L��KI�ƍ��HWn�o�U��+��r<���2,!��W:��?�~�d���d�_�jF#��C�� ��B�L�cY�,h�H�������Sɘ�paK9��J�t0��Q,O����]�B����T�|�AېQ�����Sc�)&�:(�{��M��3�!�1*Ȇ�!Z�=�hD��L��gO:���X9[�kS>�Z��XZe>�l�q�l������fR
I_��Q�,N�ș�}y�h4�27>���r�Ʃ|�i�!�Uw�o
jY�@� ��,&��+J>�{)�k�j��xH��Z�ԆN�ذ=�n��!1��˛�Ι؇WJ���ُtw�_qn~�*8X^R�='OXk�0R��>��9���L5��gr�m��d��qzϩS���5Z6�_H���Ĳ�S짙�Tu�z������`BV5�}�tsD�\���Ǩ��o�+�ygl��*�+'#���x�Ǭ��{�|zW��B�ܵ�/3��No\��8�m�\��j5cD1�����f��8y��GhPE��SǗ�Aɘ�~B��͵D��B� ��޴,� 5$&��Q�����֩Ҫ�R����/'@:T�)@N�sc��Z�Sc��-���d-�𙇘0s���c�6ɼ�WS�ސ�÷��Jaȩ�"4�����~�iT������2�G�8W��}�6\�n��}���������r�����t5�Yn���6�F����V�e�VR����`��fRh:�F���1�dxEԓ�f$3yp?kN�n���@SJs�<o���@�����u ٹd��[��WԻ�Q���T�a�P�N1:�u:��t(BT�~gkO�#~����&�2:�XF��Z�Q�����s�o<qaV��#�[�{XtT�<o]��p����⩛x�'���m��<�V�C4��e
)� Ħ��h?=���K��@�$��V��]!�������W���|(@^aR@x>�����%��񫔍�����(����{Y�AW��c��@�	�7 � ���]�a2в����k��-�N�a;����T�5'o�=�9�b�f;�קE%6Fp-��$��]��^O�=kQbֿ�S�������!F�Mû?�Q}���|*���⳨��oW^�(���I�_�w�����V��OƊ����v!�ш���U�9��n+�?���õh�vj�(��=��O_em���Gj�c��/�����܊�(5�zܨ�(�����9/A
�+&�~��w����jK��B-X��Nc��:�W��?�~��"B񄳀db.yi!��coՄ�)@�bp�ċ��ikM��&`9�
�g�͑{J^�'����GG�b+b�w��b���~?�(�E�MY���͓�lm��,������������g�n��NG����^f\���<�#��'��/���J}����礶��+��
�D�,��;qP��rُ�K��'��q�f���	�����ۭ�h�,�Tk;(J�1_��>��U�:n��K���HnH�ZIn�<y�Q Ej�(\F�_�cm��x!����1H�}�n�l�w�7\��n��;��&g������C��8-�[/R�����c\-�p�>��VW�ۡ�[)�hۙ5"�<��JRc}<�R%�B�Pb�~_I��l�Ju 7���LB��4����R�#��T��<f0(I�j�z+��Oj�)�Sm\&������ 9�a;l�H��a�h"�h�l6A�1�$�G¥h�C'�Zw�1J�/Ny�^fZ�es����Wݿ{w�Ġd^��9���ݠ2(á�����;f���Z��C���D����������a%���_M6���%�}��`ղ� *��4�ί7^Q�)j�2� &C.w9���t�F_���J�:��
����k�����bEcs^B�v
5�{<��t�mii��z���?�{�+)nF�7�o�m|T�m���^�𵝴�0�XcZnbe��Q����+D1�AMh	%�
k1���{�˨Tz���rg��<�I<*��)���*g7~�x���<L*���Z�+۔�ڤfU��vSӑ"D1iŊ��;m�3~�W�ӛ!F��~�_��}�\��j=�D����{ݪh,C��蟋]�"xx��}^��#�,�?̵GCNiI��q9QF���uy	]�i��P/55q�O���}�h^U�HXr����c;y�Ս	�4�8�Sw$a>ۂ�ɻ�b@�����?�7'3���AԴ��oǊ����r�Q3>dQ���F����T������lȘ#*z��'� +�J����y���7M�0����-�X9rĠEO�+7����$�����DE'C\ifb4�բG4�w�=}nϕB���>Մ�����^�C��[9�!943
/D�6����r�$����2c"uk�6�<}fv��	
��jX"։�Z{�=lH�9/7 �|H�E�UA��U\��� UjÃW�Ki?n��P��Z�����+f��ԆxN�K����	x/2E,���|��̉�v�о�,v��6+}Fj���4�]t�s�{u�Ǝ8�+�r��`���N4�k���(4}<~=���5k�}f20tjǓ��q�]���c�dyD�N��;r��/M�L0�}?(!`>��1j?�
̉!8/�G�p:˝o��v��U�A?�3"��x�!�(�)�ۊֶ"� ��[�0eg�_���-���R9,�"p�X� ®��͍���y����oW��؏Yڲ��?��+�5���@���;��l{�R�y���8���,@��0��@B�;-��_��b(��J�'������;�����J/�ڔ�#ϻ]�}��b�͛6������~� v���Tҗv�':/ X��֭l����;��n�1P����>PX��UMj�%lK%�%��.@�H����"ۜoDxF=��a/�
����tNT9�ݺI�E�?�t[��aɬ���R.Ʊ8��s}}���k.�>`���>wdW/��M��H�̹��V㎅�4��
	�,��Qv>j�M/������e�����ix%��uy���ǎW锂
ĸN�CD��R����{�O�P��H7=/7���O>���&�֨�+*
��{�4��iQo��b9@�4'��Z|�4{�H��iv�������A�n����>i�v�Q�y��({0��t�3B`����A��x�	�G�8��N,�$ �@Zb�!F<X^�O%���ԍ̄\�>X�����W��ʬݼ���L�u�g~k�|��3�
�S1s@h�\2?����)���cU:�^yy��lA���dV�kj��<zs����x�I���,#�@'�(�f�hF����L���p�79E��k���@���?��lF��d�z�a7^�5�F�fB�n�I+R��ҭWn����z���hi�F ����
�?�D��~.�g=����}n�ԅ�fۮ�
��)�EkN�Wo:��آ��o��ȑ���Xh?�U N�XӬ,O6c�=>�&b��,=W���{�T��#E��:��5���˰�&*�jxP��:0�g��%��2�ޗ�S3"̰�\�|���#I@m�)�;F(��83#�b��Z�-�G7aLF�XV:���)��v�ތL[�<D�c7���^����<{-�-�{����S���Ճ�@�I��sxfƘP�
�2KHmf�&u2;��)C_��-���#ݶu�o��?��Kvy�=(>Ɠ�-u 傕�]Ξr�3o4��]�hL?�n�ퟕaP?�{5�Y}�9�߲v#��/����g�٫�qO��E�x%�_Ց�����B�]Uv�����t������;3|*ŏ�樑�G��9d�O/�_��ͭ_��=�LBdd�Z�k'��9�լ�\�9�ň��w@���r�c
̙����+U����IFw��K�v�v^�����
v��5t���/~p��_j\I�75���&����`�D����2:����\8� �u8M5�nB��Ix8|�Y���P�I���ثw�d�E��E:l���Ϸ^�P^�h��φl>A�[ ˛O
Pc���0�������Wڑd[���^�ɨY�K1\�����0�Hm_;*�=��Ԉ���U�v��OO��
G��ː^9�̐\w�ۮv��y�NUp&�A����Qu���Ʒ��������UB�lK�u���#=`�#4���95��e8�|3~'v'5�x_�|)� qUv}��^��qQ/��#�je��g��ވ�@����bJ�5b_�-�FS'���3$v"Gr�nq��ה�R�����xL�*!8'��v���^��A(��'M�"y�\C�k��"��RVc�,5�x��4X�[W�^�q~j�� :�=(�nG���>ܴuu�z���l!y�lH���Gi��_ /R��*���'���uU�%�4P1��T%Tu �m���Y��73&i������<��)R�2Q>[ֲ?�W�坨��4�G�S�芖8�[ci�7�=}g�</O�Y�;7�u��U��q4�鲼���33�G������vo�8��Q}��$5|0�}�:!�G���>�lg�^<64c���A�m�)Y�	od�x�U(Tй���ѥ��䫒I�Ɗ����/w*�d(�U�~��K��>�K?)-8�Xj��P����9^���YyDsc,7GwEy�+Ɲ��9��\��� O!x�0�^�����D��@F����l�o���\�̃���6O0�F4i_:^%W��n�X�#��>9�~*SG"�XƸQ��ah�Ȅ�7G=�'7�L��9)��Ș�ЦM+G�E=��ba��Y&�mΧ��I�Lo��Z������iֻ��l�!�i:��{��$;�A��G��a�H�lMZ]	~Ӎ���bk.,%ͤ��/r>^��qܕ1�=�GW��|�B�u�n��#���zEmR%Z��B\(���rN�R�����ϗ5ͩ��_=��U�� �8�'m��h=������̫#�z���Db�D��8T rb���j�K����N?![?���b��Rh4�O?o�Tdq?�h��P(�V�ԍ����ʡ}�N�w�h0b!�>�DMG�����A2�Llc�iE�[tz׈��;��\����u���"�i<*��.j�����Բx�wV~��	���5K���x�BظG�yy�2ݨE:�'jST�H�ۃȖQ�鰶b՟o�P�,f5�:���>�n�Y���~+r]=S:����!���a���������T��F��3ٍ��g,��o*::�o�3b8�+�\�͈2���'!)嘒,op�b�	�Ǖ�O6 ������.g�Pm�*h��?~�4�y�hc׬2(T�|ҀUΗEkY-� 9���?�Ċ�[�(�1^m\ Hᮭ�cVS�oZ�~�`398�A��{�v��z�#']�8���'(a��Z�f�S�P�Tw��D/���t[��kǽ�ń4(�+4rH������j$�+UU�Zb���'m����m��)E�3_!�l&�s��=A������;��'�; $}�Z�����9C ����+�@qI�=�+u[�M�.���x�2�T�L�7�D�o������¨�^?mVW٫���(���I�$d��E�w#�k0�����Z����V�T��1?������Bڰۑ�]�!���;Z��n���������oj��+U��۠_���WPai=V=�kXDz�|��!��H��3!;�"�<�*����2H�J� ��o��w��P�~�oj�R"�֭� sj�ߧ4���?B$�?��L� Q�ո�Ο
HR�~�iu�˯^b8��S���$�+k�
43�.�6am|1�6��Dy�[�Am{�*�WF`�MT\ft1��J�!�{���	�q�i���O!K]P����4�<1Z� 	(%= ��"27�%�M�"%&�S��p������s�ܑ��1B1O-��KKTk9�~���Klc���LU!̧/Y�o�퍍�P�+��Q%#ϛ�NVU�\�pG��$4���v����r.m�f�Ԕ��[�KoO�7�U=�h��8��*J�����*�F#ga;>��x��^�Ч!1W�{'8xZ��J�g��l�tzg2�14R��(!6e*�٨w�����h����Uey�����j��3.�2GПԚ�3։/XVK'ͯZ��sٛ�l�f�k��,sE3��F����٠�|{��|�[�c��
�d��y<�pr���d.����x�|X��;��GΤ6F�v�p�,X<��l�A�5��/�/0���Yo�JWV
z��8n^�}�ǜ�ңۅ�!�z>��͸sT�y^]��j�"[2I3�䤦.Cd^��{*�lvȇ�A>�0'�=�L�>G$,�'VD����pԷ~�iT��-De�^uZ��}C�k�\��QG"͘��q�{S��5��O�h�D.s�*�n�,qI�u�&�9@�PIq���S'�l�^��`=͂�B(�Ca҂���=(?raOB�}�`��WH���Ygd�%K^��X=b�]�}�^��гzT�R��D7���M��+�O^��Z�-��h�D�uܝ�P��V��iY�� �}�e|l�U�5,����B�����$+�z��aί�I���k��{f�Y#�r�a����]��d2�$K�QR}�C���Ɯ$�ht'�g��8L�����b�J{�U����KDft=71쨵e�F�"���ԥ�{�)W-ԽS����-�P�ɼ7�Z0��XX,l�癬��}e�7��5_%��28[M�^1�H��@UU��i���2 ����21>��Ȉc����fh��)	{q̯��@�~���E�rZQ��^�Ȧ�}Y��*�v�4�����%���R�#-�I/�Q:��;�lS�n;}����%�k��W.{�c�7}?n�Z�;��'�q�N��#?�����5R��{~�~m�� k�I��[py�_�O��uK}���Qj�.t�ￗ�pZ�S���-���B��/��B��/��B��������oRRߒ� ���B������S�J��
1�.����ߌ��v���p�c�OJi���no����5Z���.5Գ(_<�>�V�xO3rc��`žK���酱��^���>��b��ӧR��㗖�II]�i1�zG�(R)��MMbo������B��/��B��nΉ
&�#K��=�I!ӛM���������Fj~~��y�*�P��V�pc��=�_d��vg��#�S���ۤj?������x�tU�[vm`�z�\�h�)^�9p������K�Z��2!y�I2�g�e%s��yL2�%ɜ/>����_|!���_|!����fCOwJ}��ڴ�e���k|+�f�z������x!c�t#������w֝mj|\�,�,��������K��PK   O��X��"�IY eY /   images/97c183e4-4c27-495c-949d-3fd800d1ff32.png��e\�-��{p[ ��[ �\	������%��,w����^������ef��7�5]]uΩ�0%i4d"d  �&+#� @�  �lD���������@��!  �J��0<1@� јUw���� �~��A�,炳�W9���O䧂;>���o�~������*�j5#O��y��Zm���|)�i��;��׷�9>�^r����y?������|�
\=����d��ִ�ԇ��Ȍ�l Ix~���6�(``i��@��e�4b�-��\�N��wBS����"D�^���_ku�a�H�c��ΟK�_�wYC�Ѻp���8��& I���5�aǵ{�޴���b��l�/����䍚Ԋ��ޒ�aÖ�¨�w��Ce�R���r�AüE�Wq�������D�L�����mImkI���w����c�}m��à��r��?�;�{~��IRB�'uϔ��4�7��M��+G箷d^&Y;����_&C�'�Vk�4�f��o[q�(E�����5j#��a���ލoI�����jȓJ�	W���k���$F��v�մ���5R魍�˝�\�M�N��VK��+�>��18���Uw�۵�d�f�O�_���<.��k˭G��9�[���w�U�4�ԲM�py��A}�U
?xP��rP�(;p�-J#��銖 �ixLD#=A3~�|C4���j�*!Ǆ#��y���7��v�K�#��G��\���� �4���B�8�A,����R��@�	�<Sj���qW�|���)6��
G�fW�&gL���-/��-M�D4���"�(��@�u�hD#B,�2��F~�-Mo��×}j���n�e��F�
9�y��rPL�"@�*4vO����1�̲)��;9v<��s%�M�|�.�.f�*b��j3���al͋�58�Խh���L.���*�����Q9�S������-�l�t���D��6���.�A,6�����z�_X >j!B��!�Vxܛ�&A��V�ˋ�*V��~U��G��1q��9l�Q�"6.��Xg��_��;�6Ԛ|Jȉ��m�ұ��;�N^?<n�>��&sb���-�����������Iչ?S�=]�V�y�w6�ԍ��(e�d���`��6^%Wo(�]���k�V�E�����E����ңm?��-û#\ٸ �>�}�����q�����/}WxA>ҏQ�~���$9v7��4����D�h{{P�%v�ۿ������o�-k�_�8����<f�h����̶�(}܁ ��$-��#�S/�.w\�way��O�^��Bl���[O=N]��c��?��H�`GͿ�����d�b_m����J3�V�_����1O�%���O��:]>kj����)��	6� 9��h�~�,�~���Խ�q��|m�̙='�T?�-"����dV�-��M�G��,�'�8׊<
-����^�%�	<�V����J��׿�gO������������/r��[U����8�$�cLf{�兒���_$]G@�H:�Gm5\ݜ���
�&*9Ǿݟ��r6�rKu�TNڤ�>�%����jA�\:�������R��Ф�|F��ᝥtx�G0fAo 8�M�����僰_�F��s_�b�Q.�'X-��
������/����E&�,�;��ʀ|����S�ѹٗm��&�I��d�kE{ι%�����*S�|��: �a��O@I�s�s��Sҵv�j��b����O縉�s�\�z���C[�%׊���kL�����������|�%����B��O���d���˰d4�:���⢎R�e�������.�[A"���e��?
��
L��Z�?�{8�����l��%��R<e-�Bu�0���z`~�]b^�E�����vhE��{9�m��y�nϩ%�-���N��y�}C���&�T��ӍBw�*��ȇ�`2�6&H�+Z� y�á����y�"^��e_z����s*k͖��U�5����G'4�NP���L�;�����<֯o������q��W�"Գ�l`O`�G��q�b.����9b�K�zx�]��r��a�V��}Z�z�Զ�ZC_$����f6n�GZa:�9jQ�	�$[�GE}��[�������� f��MRӃ_c?��y`�C� ���/�3�2eg'�Z^���mob�xH��E�WD��3Y��y'�l$1�Z�h�m�4F3G��RQ���OO��u���Y��n/Pl��A�X_H�]�m�����>��?��/@����Z-3P�%�̯uRk�T�H�����P8y`���Ca�[�ZP^~TJ궴�Ǥ}aY��D<o�H���t�nr#1�Q���'�q FRۍ���QX}.>'�g��R��h�)�-^�739��'6_M��
����tjez��`ԡQc 
H)Ň`�k�<�� a��On�D�,������o�^܊8�㈃�#��b��a�k@cї����S������]ZQ�qYڬ�h�u��|�}�~�@[��}iފ,���V�q<�D9L�B�y��D`�#:j�͊�@0���m�ș�.��K�����z1���� z�m��n�b��\�� !_P���aM�)6�!X�pJ�.����{��3n���/ʲE�J�Y��W�_�L�d�h��,O����=��@E��2��h�2{��AקL��V��bf�Z�?��Y�����\�;;J�lw�\�<\ќ�L�+z���0 َ��)��$�S?�n`��lW��m��M���@�g�����f��o;J�6��������5X��뻈���t{�v�p�B��Ll��+7lkD�\O.E?�6��|�a5�dZK������]��@}���EI��/�9qk��N@o�Y$
es��I�+F�����U4K��-	��c�w���~�X�����cM��:��ή
v^>�j"��<�Y:�������l��5,cf-`b��ǭԯk����)ÎM�dZ�F*-{�X@ɹ�Vju�Gg��"˓DU��W�0����k���Y���.������Be�����?:T�O�VI���OOO��������U��.�W�q//
�uu��WTD�t�S�	�����|�eH�s-����/�4��ٽ�V�y����6��c����e�&qt]���xy�%yZN����S��`ՙRC�O�ޟ�ó�C�3���ܾ�Z�Vepۢ�q�"��<RYnUt�ν�v7��u�x.����m�Ε����W;�Ț\���%L�����몫I��z�"�ك�77��(F04p}��Z���}?�ՖX�d��mɉ�*�:�����*�:leאs	�up�5����R��/q��WZ�&��^�\SYUQ!S�h۩SRe=�ۣ�޿���Ȱg��Fۻ�~���l����T��.�5���̧M�v�msZc���7ww�G�Xb�J�r�G��IwK��l �Ӯ�3��('c��F�Q<��(^�ۣ��y��Fk�U�۔�jy�� �X�^��xb���h��"�|������b���9�s����n�fT~yu�U)��5�?(�\}�����RÞo�#m\T����c2�ƟN]ݱC�	��Y7������y������� �
S��RL0
TL!>��6�ɱ�0w�J@l3�in�u>U�4	�A"rwʗ�	�P���ԙ-d��T��/��$|��	��k_>0����_��'�u�'�ؐaZ
Y�ۧ{�3�f��O�M,�k�����8??��Uk����~�gd<z�,E�:�Z������~kV�����%�k�>[��F���¶09JS�@��&W��A����x�2��=z���8�*��8<�Z����7�C��J��%oE0$v!?N�܆���"DtxVw�t��V\�~�z�׿u�����+6|��=Zq��P^\K����>30Q
��F��ۭ��7�I���da-:VG��e-�˒�kv��,��B���}	<�'m�`������)�땏�y^}�:�i�>��?���Z���w�'��#�T7��tT.'�m�O�i������~�Ͽ���ۧ�~ ��2���b �E4��?ؤ���[$�>��#|�d C�w��P K�$��*�s��7�	�._�®��:�0Q�8ax����D�j�*T������!�Ժ��������6�]EE{W���mH��Q 8��F;!�V
�dv�?U��T(�����z���:��3B�d�G5�==I���7j��zK����/�p[��uJj�z��^��d��XdRe�m���J@��a$�7b.�ϑ�!��%/W`Nd��B~]Vշȹp `�����~�`"���)�_O���MF肠�,k�h�a��x`������N�"�+�bΩ
pQ�KR<բ�<��o/��SF���J�X��4-ɍ[�{��A�]?V�0���H����i�4��|����)pY��Q�"703~��\>�/�\NI`d=oa�-OO�F8��t��D�9�<�'S��܆��8y��=�=f�#hy�|M�뮁��k���R�VL7���`lM���}2��!=�n�?��ΜH�繁���2uf�o����$��/eJ�n�!z,v�G0nok� $�ew�c�5#���ikˉ���Ŵ-3I�ihR�h릢Q���%�3`"�B�DD[������a�|T�%r������+W��Wօc@�����8z�N�G��G�**ܡ��.�'��-ϛ�(���d���
�Oo�0�����k��+��8*��e4��nZ	r��a-�T��������{?��z�o�a!��sB`+�|�Z�pů��r�1(*�2n���N�}�W������_�R�q,V���,�R���ItzȠ���]��0Y�*S���hBw�/��|�*sn����y�C����B:�Ym.Ϣ��o�!
MLA鉨�CՆ�L�� X��pۚ �F`�w��06������_�Z:FI�Y謨v�_Y�c��n1��ϡб}b�GĴQ[��~����^���)S����|��/:������q]:� 7*eFD���������<�r
�����v��u[=]hu>X�]i��[���R�q�z�C�����l�����J�<v9��h���@��q��r:���'0mN��ʯq���أL�K��Y)09&G��wd��8�Uw늳0��!bC����)BT+|��u);[�j��1`� ��&tNW�I��62΀��@WEV܈'�d:�b�xּS�$`y�������B�QBj���J�Ť�T�Ч>A}��Ak��>����7,,h£CIg��	���³_��R�06���"�WO�"Ʉ' �$A}��	���\�p��[o	deeƫ�<	W`���##FDM����C���ȏ������wS��s}��Y���z�7��i6g&AYd�	l;�����S)���_��2Ca@��O�Y?���ɸ��ƫ��r��+�)�|��m�~��JG���Ƴ#8�c�{F��h�rܯ��c8�#�k挒�t��$0b\�@�v�����8
.݃�Xwā$��ǋϵ�3�.�L�3�|���]\h���C�(9@�N��n��q��X=d��&�;:��F�V1��u��,��rB�/1�t߾wm����U�(�}��$-坴�jw�pk�Q�J��jl�o��Viяk��$Fxm�M�]�H������r�}Y��oP�G���
��iEjof��'U���[����6¤
ڻ/ (.���W�0X��x����4�	$�IH0��o:Deკ�t��u��%�o+�ԣf��d�(���X+�ˤ��~�<�n�q$?���|��(��^s����Ӳ^�}��o�=��^5v>A�t���F� ���EC� R	���+SZ�"��+�_H�%͢g�@Y�����G�:5�g9�:���k@k��G�:K��.檡��'p���(�pj38辕��J��o�+������������>8�: ���n��=��<�O]�L��}��i0��`~��7���؞�/����چxp�?Zਔ:���� ih+��0I��R@��5K������yɪ]{�3<�f�:KN-s�U������5�r�P���'��ŸhK�i�x�ҹd�>���U�R�g�1�qۦ�i���s����P=�e���c�V�kO�읤FU�w�@�Cڂ�;���!��> ��P��'�"��I�@�<3�JyJ�Q0e!�3��$HD�$L�� ����Y�����(a1���;�Yn�&�A<��^?��]ݦ��,��L=�5�|9ЂOS�#L~АQ%��~-d������C��5F80�`���a끏��핎�W �R�v;��n�^EN�s���Z�����l"L9�9 �,��cWrw]�yk��i���27/��{�H�s�ְ��8_��
1�?+>�Xu����A{s\<��m�|RJShQ2����<ؾ4���
�7A�
���Q���A�YX�P5��Q8���/@Ze___Q&Ǿ��R�C^���RU}�]I�o~ïUC8�p[��"��Rə��N��;8І�郋�,��Sռ{�,��^_D-��$�FU��2�>�����UQ$x�]@�Դ��V��v��bU��#O2�o�����?�j���Q�.$C��l�u��c��7e�|�9�:ϯK���S���AY��
a ȧ�k�Q,c���^�_6��D�����D�f���UPqX`!��1��!jF��yd�T�>�������l1�xy~�~�ە��.�."!��A�ޮ�5�pG�ؒc�7&<��1v���#�4˳�����~_��!��������U@��yT���c��K��,�s� �|�0�{���ֺ���~B?[ȬiS��cҾ��{���� ���75#Ŕ�Ւ�h��HOq8ڴ�Y���5�5?A��xS+�5�1��<���9�O�gW����r]'E#x���c͡a֨����Y��E$�;L��e����eꙛ|��L�p�/���F�Ij��ڝY����d���(>ٖ�����(���3�?C��?cr�2p��H�m.v_���7�y.[w�����˺���gw4�u��������W�a�Tq~�`���y�%�0��	l��5d�����Ǆv�/�f+,�>vf�i�BW�!�Φ��V����@pK����a����P���(�h�c��,��A�L�)�mε��<nKU��>��訍�(�3�=Dp��Z�F����z>K��0�Ц��L ��Q���-WCug�B�y ��rt��j�bmqh�#��U�h�*�oo7�������mΣ�G��qJ�u:�N��v�L2��	6{���il���:�t�?�c&LS�
#(���9�׮:R+�j� "푯��&s��2�O{#�}g
e�|�36^�ls��ը6&Xk��"[��Ğ�]@��C_(��M!#l���L:N:��I�զv+��9sSMwޮJ>�k@�"4nE����]���4�f�Z�&og~����;��!J�W�خ�|��[��@ ����+F�����nJ��`�<�a�rm�3 ��J�ޮ��>J
��)$y�a�ǩ�s����ؤѭ_�Y׼ţ��b����S�VMlU��ʲֳ#Y��|�$�d�n��bj>�VS��K� #�?����%N��+�����)V+$�R�5������]�������,�W{������G�"��u~�����5��*񐲡���=b��j;N�:�#$	��֋�G��!!�9�Z�Y n�`ic$�r�܉��p�D���(������G|�6�KJI��edI�^A�4�|�i2������jI6��;���c4z�3>Q��+s�/��Q>�a]����T��FT��+$���F����&m�1�U���ٯ^g����Tc0s.�۹[���X���}[̹�@=�/�^L�.�sW� q� ���6�2�P b�|�������`����{�j��2L����T1���c��ߞ"��n��}��,��Q�b����UC�A���z�H� ֊����me#��	����P�Χ��E���
��A��t6e\L��h��:h�Ԅ�P���N 	�$��#z(�m,X��ͤ��J����x>�
%���K1z�H����~`1����=�Kȼ?����?-r"��x���En���8'EG�Z�������{�K,�6����aƨ���3ڥ���6~�����T��rT1
s���l��6)��I�q,���*Ċ�WZ�$����~�T@�ڷTs���~�X�k+���`S4�kϚo #I;r�iV�~ޕa�����
FàG�c_\j��F�!�_�Wt�U�1��c�?����KZ��ᴦ�u�p�9�r�f}/��d�3�$����J%����e�+��?tE��V膇����x�a �@*ꈌ�R^C��ݖ���h�։u�����;��c
]5ARD@!��<����u��<Py�m�u�ά@,a�X9�7�������w�E�?��xf�\��1?��vX�P�V=�K�܍�kN���Ӄ0���L��.�1j"���lvJc˖�"�%X�>�~;3�f>��.�+��Q��5���u�h�ӷ���PL��g\F�L�e�Q#'}�界ru��X�jn�Tac=hw�o��g�Ii�
ì�L���ўK0�$@o�������X�#�K
����e���C�B�=�H�M�ύ~A���ym�b0o��*�i�(�K�1ӊ��������U�/~ͼ8�/�?ԓv��Rם�u���w!O��*ΝM��p��⭮�靔���?�Iq��N��\Mŧ������6�O��q�a������`�|��:��tVi@�+�HI �s�)�˘F�{2
$�lE��Q1�\\}�e[ۢsv�N�ug,��(�T��
�i�ޯ��Z8"���G�9�������m� ���-�g����llV>��U��E��x4����Aq37��D~P�پc��^��v�֦�\��u�`"�>�Ľ67�o	�j>��t�[0⃡�d����8'_F2���*o��B'��npX���eٝ���|b���l�7O����ҰY��3���e\����aԗ��<' �}�$>�9�Ͱ�����Ԍ��FDD.I���jo���B`�ˁ!|������^F/#`O��.f�LCwr��t�#�Ӄ���O���Yq�vK�crI��}���l�:���NEv6�,M�ǻ���*��fb}�0L����V�	^���yu�&���g�!����������$	��Ws��|�Q��|���p��[E�@X����?6�c��3����Z�������nO�/4w�$.�d��ג�p�9�⩛5�"�4apo�ఔ`�	4�cJm���?==�(��%R��ҾO���k� w$n{^�H��c�R}�Ȅy�9�5��j�UBs'/Čb�\-}��|���ً�*Ϛڱ�y
8�06��,;�EW���d�[�~�����.����b��^��b��{�;�X9���d;ޝ�V#�(���UxF�C�N�ǂH��ʵ�o����\���2+��ջj����|�닞¬Ь#�D6<��i����b�ϋ��e~fWsQ��K��\3KK�j��m�04�H�	���].U�v�m_��JK����b9#dPi��9CԴ�^_E��Q�ժ^���tdG�w�hp]��bs�lѦBU��)��>�C:��U�;Ξ�YWw���گC�phёO�ˋ�~�(+O"���誫�|�!�+�p��y�GyT��/����^u�l���l8��Q�˓������{�C��\$�M����`,3l���	��Ήv�엻m��P��KE��*�h�*���`�����(j��)(�kK��kMc�-�<�_�c����F�e�-�;�E��N��Hٷ�#K./����7�����!g� T豟��]�4���m.���%������֐}/���=��*Y~q�<�Xu���gE�Bu���(C���Y+!o��������sSz���+��a��ٲx;,�@3G�r��^{\u7��n�4��""X����V�pd3Ič�!r0p�+S�綘�<'w�7/RP�St#9(^XX�8�7��b��k��naZ���^�ZKa�
�hhEA����'����J��`pB;�B�\FY@�����翄c��s�۔ظ�p1����Y�&�o]\��h�6K_�S&ĸ����Þ�� �xqE��z���l>mҵ��q����P�������+++�J��7��ө�j�}-,n4~k��N�m�d[cC���3>U����Ku�]����L ���h�\���jݾ��i�E�+�6�7�dH�=���#tJϽ4�yL,X�N��|�K0a�1)F��ql���M#Q�YhsԨbkC�F����t�W�l~�UM뺡�f������F���ea�m�Ŕ(�F�g�]�7F[q`(5%b�]0Ůu�C���At}��Ԅ�BмM `$���O,��R�n��)<��F�^��1BWC���'���v�Ĳ/�W[��~k�ʬ9�Ԯp��3e)-%�Uh">�]�!���|e�J/w�`��%��*��p���g>�j;�!%M)̄uh#3ޡT��1VF}�ko�@��-���w��w�$�d�|�xS۾Z�QJ�B2�0P_�`�U����g�Np�����7b��7��y]#���/�4wޭ%�(�_O6�rs�Fr�o�ttN|�%�f�קb-#_��r�����%.��r��Mg�~�G8��)�ܒR��V1��{cҤ$�\G��ߛt��رg����f��%R��*J�[�fY�i�`�A3ԤN�f�
k���N7�ߣ�@�]&�-�^ɮ����^�ֲO(/��	���"�%��y�:�6����C�v+��k�wȴ�3��iM�������b��S�*���*<�j��b��V[\\��-������#[k�o�$%�@�����;�Y���ş��N�Yd��/��l��@�@��ގ0N�>3̻@m�ņ!����]�֐9C����B�P�7��C)�+��&��p�l=�\��:B��p��/�|���[_l]{6��L�B�C����W���?0�eWz�\t��8�/]�eC�t$Y�cz�����D���7sUo��|��:�2��@2��������wל@�1'ܯ$lK�����4�$`ocߌ�!6�di����"�E,C��s����^�@�;�m=�~b9��3�w�i�)m�#3�Nu@�����u@N��V�KcO{��+�<��#|�p��ܱm�%�~�Q��.9ܑE{=ɽvq��4��ց�#�P�X����vaF�u8�����J;�Mk{YDȕ�{��P�JC���L SX0�P��`�����G\4.���A��U)7(�9c~Vy5�h�4�+�'��M9ZWz��Ԍ���A_�����*�6�a�$Jj�� ߘv��.�����`]�Ѐ<k�J�������V@v8��X�c9���`M'���A=��ں`BKH�e/`�d�]0k�����S�hZr���`�����R%ȁg���B��Tl�$n�������K�@�rߍ�n�Y�����ɶ0�LA�I~pe^�Bw�I�ZG'�'�0H0��:�N5�u�Jh	�Ĩ��5�c3���M��lL��=�[�MY`�����q���gDu��p�A1��:S��2�|"z�4ݦ���ɘ/��,�Ҩ4�%t���S�$�LO�Q>B3�NL��2_;U����=7֞������&/���i9U�a�x������"8�Foc�caEޠ�i�
X�a�v�x�]����O�5g~1�i�+�zk����FD��r�qD����p3���i^��N����� �����&�S��[n�S5�H�5ĒJ;+�"� ��g�����B��荋x�?��J�bC׋P�+�o�#c]!n"\
Kɚ�T�
�6�i�3��p�\}�פ�a���O��Ltg�D���-ͨ��w�,���2�W���P~j��$�N�vsu�PpN▹�PO-l(G�Ƿ��r��mQf�a�=]C��_$4&1�� �Dܨ�(qqѸ~�)��:0���E$��ZK�����|LL�}&@ս<?����+���?��A�|
Ke�):�O�c7_ ƹ�x;��4�� �BĞ�t��?���]M]�����/ bs��O8�����5�P���J��GnifY!���j!&"zr�&�5�<=�Ԃ�
�ISx������pa&�G������
uGG��	Zv�����ȳ�*�^��RB�Z�.�j�D��f�n	F!1�֝�3e���@VK�Dێ�Bl �@��^h�ց	��fw�bJ�4.��晌p����ٷr4jm�{��('�'�7���@��G°��Z��q+ip����%����Lm^� 1��ZDQO$"/���(΂��j�.d%@�aW���8��Y��v.��Kc�����>.�g�ܐ=�ְ�����&��5\k�
��}^�szB�9�P�UK��t4�s�����c8xg���RX̰�3X~���o�\[��ԶT�v����y�t�y��;�5�1b(G(�mB��K�7x�c/�X����ʎUP�++%l�|�NҨH8َ/Aǫ��~��e��H�,�A�׽�i�#J1�C$2�,$+�Q�@������T':V����$R�tZ����yђ,���Ԟԟ���|�c������'���F�{�wk���7�#�5 ���Gb3����i�DbwG��v_��~FI��TlߜA#�`ґ	��A�IҎ�3���O(��]'!p���g� "U�`1\�P��eu�	m�F�~�ʨ�;Z��vDG��B�޳"�ˀ ����E��4�_��U1�o~��65���{u�E��]�8�HD~��<�����oGycm�2�?9�!B�k����%6�,,h���8�?L�ZB9��ؽ�z�I����|0�j~��ށ:�TjR2ѽwR ��(��bր6�X��TD^;�Q S�V�i�V���~��l	�C�@�>~��Ȁ�қ�uDo:M��V��+�SKL��a��l�hQ9狅<��x�)8��d3�XXrhY�G���%��[֢�G�F���"�t�ON��)�S�5sX��db컗�������|��ɔ�����59�ސ�b�HJ�4�*Ej<���r��:���:��Vr�)F~i��q\u�F+��s�_�/�rN��U���K2'��2��������.�N�"���;��U�
%��T��v,�}�i&)n[�o7%��2A����r���#�P#���}h��4�%���'��P)��)p��@�Ts#�^8�st^��Z�����)�CE_u�J��E?�+cDTJc�QO4
�-����w��,T�2�;��R<���;W��/o����"�e��Ʉ?=t� '�SH:�O1��pjK��L��P�ۣ	eCI2�2��w�$�6â�T�H�cB��O�j���X�>���S����f0���sh���7���	��;���(5���?���/���3�ny��_σ,��4��
���׻eN)��3�6����n��ARw�����H�I�w� V?�4qJGI���SZ�T���������m�O�J����W{���<�+�<�C�?t�Z�AIA�3� 6�����PRb��C��j�W3� կ"a[}�lLKl75�'?��Y��u7w���;�}m��fy_��i�P��3AwH��/��Fw����18��C/zyX�u� � ��c�@���¼�E��ge_)�5���>�@ �a�%?��<��!�8	ikcc�Ņ�_Z�V*���:c��@�އ�4�A�D��%-!U`G	Zw���Y�I����8Y���3���p���!�,�T��獛�>�z�R��0��D���FN�����l>GJ�_��?�n
�kY
�5��|O-)~���!�7}C��HD��0��q1>��I�+�!�Yl����,���LMƭ��8�Bq�Lxb�L����]ꐕφ���|q��'��S{�c�P�׿�����EEu���8v�z�Ν�9�����Lς�_����ȝ7W(nC�z�����.�� �8l`
����yw�4�2k�P�NQQq,��
�����#-G����� �[�3���\�Ԋ�/2����c��gp�>�V����]@�
A�#A	�����^g�Y�-���F�Ʒ���GrlyC�!6���U_��`���Mafm:3��*o�܁����v��q8�����yVV35�}}��Wڢ]���S�����P�x0
r����~�ҍٔ���+� `K=�x�[p���Bz]�x�@�d�V �! �M�	��X���n͈i���A���E6�-�a"pH���cGB���1���L (�@
DS�.��t�Bt��5u������h�ll@z��;�h�����d�Z�_Ƅ��0�t��?ȁIWQ0�l�a�J���.�*�%���Hl0q���
�����!�Uua��S\��сDJ�����	?�&
a��t��n�No�y�<"$) �&��~	�.�ͧ:�	�f,�]�旇�Ů;�豶���z˸O�*���EG���?m����Pb���ƣz��<�� w=�BҒڀj��c#u{H�
��K��(Ky�)�6{(ߖl6dO1K(���d6f�|�>��r�e� ���B�}��4&��ڃ�4X[o1�w��g�.�A-�0Lh���<�*��4,"�y���'Ii1���-��蚶1�����F���]���I�W�]|E�0�{�dM��ᶡ6�������������~�$d0�����D8W"%b��[�R���3��|�ؽ�IM�6� Ɂ����aۼH�Ze�ؾ#.N�����f�@���r��s�
�hd(����Io�j<���zH֛�z@�ɩ����_�uE*�'�V�ap����h��;�~c�(���!�M)Oi�)gt�]Lxg��	���#��g�0��B��v@*f���0�,  �K���J{9J��p;��ì	�_�y#�@*���~�i]s4���Eh�����z���{��'��ݗ�����J �s�+�����$\sR���*���p������Y�0���d�,>��i����~�ڼ�'��=��0R��1�,��I`'�#f�`��CUj�S^���D�;M$4}���y�<��0�48����L���M�qb�����BJAQ[���a�4T�h@���e����Y嗄�J{��+�i9�%�ǢϺ_R>c�A�$ @�P0A�#�����s���vr6l�HPFP�i�2̸`�@�I:F�-J]-8�^�h�?a1�n�)�fX)
��5�y��UD�t��@< t��e�悙�/��n��i���@����������i��ԡl �?��BZ�mB���v�~xMDے�3|Є��;S���`���	�z>Ø��KK�ٲr�'Y�k�[`!t�ųK�P<��zK��:m㞛�0@���EMN?$����}�A(�V�����F��C�I"���BC{��$R��KQ�$�?��?�N|����xC=���ql���F�]f�tK������ֿE�9ת�Ϝ��T�i[Ռ�����|��٨gU��+��@ZV���Ģ֧�LN�fY��'�sSvmZ�q���Zҍ��!mx�w�!0���3�DGr�(d��(q[��,�ַ�Cd �2%�p�A���\5H���ZY1�l���Xڌ*t�*��;<��SH�j<�+o}���Mk�ە�1�N���xe�G%t�kk"�ՀSr��y�B�kίt�_$��oZ�T���2eG3X)~������84FL�k��o�-��wI5�d2��jB�g� j)����/"�kS�8	�UА�kbZ�K6D�ǏZu�H�\�hc�ɶ�8�p�}��G|)d�t*Ȝ�=q�'�yy�0��t��
�p��*�)A,�E!)�[�w@Bay^����$��we8V����B�\-� r��,!��>cH8M��o�)�*�4���8UJ���"����>���������`*��p��{�n�h]Fg��0T�3d�f[r�*"��.�r_���iF<�̼3����ƆN�p�������N9ݸ��ք�nI�2h����&~7�~�e)Q'�����{�Z�a.J}WʉB9���N�-��v��of��.�\���U6L�=�Y@�7�	杀�s�Uw6-ƽ%�4���@t���� �t���v`����A����h;X� '�,�B�E_���+iC�� Q֖-[�q"���f�w�}7�ꭈ���]zŒ�+
�3�Z0��c�m���)�!�2)jUs�>zu�˴j�f������B��*�'�d��� ���B�n"ɚE�=��ә�/]��c�/��b^#m��<4@Xw����X�,���*E���v¥tՁρ��'��`��e���[�lP�����h�޸� ��6@���qV�KX	j�����p"I����]��oo�9K�n���҇�p�g�r��C sbvG������h� k l�"�J��o����"���z�N1(��g?�g��فo�n钥�Ϙ1���-�Od�@��}�m�N��a�9�DGqgQ{��g8�/q�ೞ�Lt�=��eˠ����y9�H���̝;�Se"���{.� @C���+3���Id�Jh¢/sSv}����8��4��+���� �C�âYn�?��]���X"�$*"�� ��c��At�_;���* �&v*GG��L�P�&Gl�Xad���^����_� ��!C����f���������d`��X�^�#�Iރr {B���7�#m	�Z~�u���(�Ţ�@ =fi"���K����ԔT:� l��_�}���~�#,G@@���`1��*2��5��P _��H U�.p��1DO��'>A31�3v���B\_"���9܏�2��rHY��p9@��\記YAzB[@�]��tNY]��㡝���@��"3$ee�r�p%�D#�L�P�=��,G �����Ѹo���� ��� Z�'�p���>e���.��#���o��wQ?�I��aQ�,�A�(��K������Da�N!k.���������*΄k����Q%�����'��\O�>���4��;DlLD�C�d�PD�����
d���0�E�
Tc* �y#F=LM�^R��K�!t����ߩU^8�_���ԡ����ld;8��\>���%�\�!CX*�����}��%K���mRd�9��) 3�E|�S����v�1��M�N;���c��Vr�UU�q��X,�5���;bW�Ry�GÇ��XĦ��ZY�p��/D�\�n���|�v�,�3X���e¨�,�3�=H�'�fx�,���5D6�mao��F��xa�1�	x�&˜���%U%�@�8� g J����T ��~ɒ%�DnP�)h8�ԝC����TO�>��< � b +��#@�
"
�a!0���`�0��V}z �Tp>K�K�'��e|�녕��(���'��@���_�2;D���_���R�B�B�<����z4ˠn`�f��lS)��^ �x����\���� ə��y��S��0��<��nm#��`�g��r�,[�凫Yjǖ#`GHP.�.fݲ�	��N����-ā+�D��, ?p�a93��s�B$S�/�؆t� o\C4gd��k�Zok��40av�%�y�V�!�l�Lp���P�9��	���'�S�0D��Y��\���7�'(+�D��C&\N߶���YйY�i�$�Ơ��^��e�{Ǉ��$�Ph��b t��:t]]��t�eG�[��ާ�XE_q]$ٲ�g����6�+���>�H����O���d2"ݫ\&,˖/��"����&��>ș���(	Y����I��y�x%۱	pd�W��C�Ůz����f��ZZZ�U\�hغd�H��I����Y�P�*B[;��0�3AR�Ĩ� !��tS�o�ы!�x���YY'M Y�3*SOa��T����5ϰ�\�g%�@Xr�~�_�A���$��`��uG�����>g���*�L0d?�]7�0���`��o��rx��͡T:N;��T"�æt�#�Y���#��K��]�i�0�> [w��e|q�-9" ��p,�?(��^@%O��6���r��cP�h��%p
3v����I�Eڧ�ƀ	?���rn�AxX��R��јͫ|ȵ����8!vLX"$� F,�	�a��sNd97�w[�P¸zܱhi�����0�$�A���=���mu��5�\���!RF�@tJL+1E��/t8	���<W��\=��l2<8�l������C��R"�A5�1���7�ܴq+�{]��j +�D��^��v�A�|-&%S��{i�^�s?{�u�ԒR"%G��GV��Yl*� ��ñ��U.��LGw��;y���`�K"/q��;!�%�j� �=|���`-��6ᆭ�~��`�X1��fN��]�og\=c:� �taǨ n�Gc]L��ٌX:*�?��;CdU6C�u�P���U�r�0�10"#���zv�bօxqL)!Q@'�|"��s�� �@���A�lbׅ$Y�C��9���h��u��h�ȱԶ����p��jK�l+F�T�b1�J��uS]}Ŧ��9��Z�#5�x�J02���1���3�z/��+�T�!2c��U�F��p��X�N��	~H�S�9�1r� �����B$�,۶��dɒs*΄�un�d,�H&�,G�1T��e���,�+��l]W��eDp��	�ʻ[��u�2V,���2��v�J�V��<���s���:��О�1 #h^��Ndv%��ۯ,��)�) a���L0�%R�t����9��葿���珔L�����*��cQuM�z{6Pu�G��z���C(ѓ�_��z��)�Ĕ��L��uc2Dď�U�����aܕ�`�~�w�ل��	�$4ъe���
ڣ8NESFy:�	��H0a˲lii9�� �sЄe�\Ĭ�c�;N���=�~C��
��8.���d�:�fK0����G/`L�WʔN���!j�,��rv�֡i���Rs��<{�ˬ �UO���"4�B����5�j�אَA��ɁT���>���2S»�1�.��:���9��mS7]��[����J�]1�u��^&��&Ǎ�at�QG͢�.?���g<|���t٥Ki����%��5̂�b� <��S]����aѢ@�\E��6+��ܩ/�2(69^pI�7i���l�I�H��1:f	��94 �V�q�����2�z��{���%2�	x
��ߗ��) ,[���6)�(z��ש������ib�U�4ȕ�`�|���.��v:7Tv�Q���\�$SNc����k�ԇW����g¶��pH=Df͘�}�������"v����?�-]s�w�Pu�Jۈ��{��ldQr���I�g>�x�}�Ewu�袋��G}���*r=�c��k,J$�X��\YP��d�:���-s?F�%�q�m�䵰L�0a/�����#����I����t�@'f:��g�l9R��e�축M���qKȂeY�x�p!���B�uM&�u �6�_#��} ��ʕ�Qo'Bf����=�Q,�_i�r&#)����B��v�w�E����g����R���5�G�̚ <�H���{�5��X�%:`�T�x�G_��{tǏ~C�UM����2c̮���6-���L�5)�s�1�ŋ΢Q��y]��6:����Օ�ɠ:R^�#"��lJ�:��[p(��_1������:�LT�U�~�1��YO��@X>}�\,�N��H��8儹��>;�{ ���/^|vESY"w��0{��ݖ� ��;�@��]�{[0�� ��gJ������Jf�1И�V��#��Y@c���Y�0!�	�����~���e����2�DF��ش�t�Q�i���я?���wQ�WQڱ�@�Z9@��z=�϶�]<����(}���c��x<A���~�ӟ�A�=Y��p�CZt�-�y����g* (���
fFy (H�3�~ f����'�}�, ,�$�o1=#Ć��f�2��R��yB:���+V�8g���{��{ʐ�|#�e��[%�/�T�NF��Jv��F*��a
MES�Ҏ��Q �W����Lt$A��N^�������X�Ɯ��}�Di7����lJ���o��1C�l#�d$)Z�rV��fq��$UW5Q�!rU�s:}��̣����j��t���"��ck�{��0�V�����+G9�g�Ad������* ,�vp��������a�f��'�E$	;��q:���H�l��� �ͪ�m2��
�n����Tt�� ��	O&�°��̒�d�w	�ֽ���v�L�C�꥕+_���8Y`% 1�,8�����<��������_C���҅��4t�8:�������(ք���jiJ�{��;� �I���y����$�4�B�
��;m��! ���]�E� ��C��R2��H,ʻ��%ۈP:��6�Mv����7KLK|b��>�zM�x������;Fk�;�d���S�r������W^ynEA��7j_wkM�{��ә���+�k��#t�~� ���5�	��p�Au���/Ȏ�i<� c�x*�dv�:�7TQ�LJ_-���1�c�Ow��|�^x��`��SQ<��a�r�}@�1�2Ps�4��v��C��I���"� ��ҞK�!�b�h���`��b�����qd9�0�8���L����e�BLX|Stv[�g�.e�\	]�5
�lXo,�dS'�Ax��˖-;w��魃id7�l��zk��5)WtxBu�蚯1��M��5���ܱ�L�|�U��a�r�,���o��+�tI�h�.�a������������
u��N������c1*Ή{�巍~P�m�
��Kv/��f6��������X�gY1�OCԂ5)����Nd������M������0_t �2扦��]a����ئ�{���yf:�f��0a=�ד��L�	���g�BW�w |߲e��ms��Bn�	���N��BŰrl@��)4-�A�s�lp�Ż���� ����~4d���ӊ`�r^�����TXm�r��^87{:�w����6�p�	 �~���ֶ���@��ة�8]�gb`��5�6��$"˦X,B���c>��
̖#5�\_�,$G�kC a>L��$yn��qҰ���Vˢ���F�r�9+d��%s<��[����z��dG� ��,Y�+�rQ`�����I�2��\�U�aܷ|���*�[Zo�IuMB��D<E�U���dG���rF2L9��	�e��$UF�4�lBJ8$F�)�>�隱x�рa(�=�~���2U	kʌȈ���#�wf?�	���ʡd*NQ+ʫ9~ҴȴmjVG�M1\^��0_������`��{$���З,�o[#nu�Y�A��+�-^�'Y��%xj8�1(+���[�`Ov�0�o}�^la�Ul��>#	�		��|�6�%׍S�mQ$bR:��^�8���f�u��B�j^y��yWt7�I���ό��"�r= K��VObf�|��ÑL��,�@�� �x��">�qQV^�~������G��xG��>;g���)��m��.^����3g�L��/G|���M[Zo�%:&!cF��H-�`}M��{:9���C*K ��X�1x8�I<DT@e��ȳ�>�ɑ%яhf"����908�(�
�8O O@X���Y�Z7����]���R*N6�$�IɄK��"v��$�	"�!;
	1j&)ׯ���GG��<����;63ʹɧ���{aq�	 �^�&,;x� ��b�Z�[3�
�w7�zup�{�I�`��L�ӎ�d�d" $n��V��Ӧ��CS�΢�j��E�[�|v�T�([v�f���|���g�������I��?��o�C������f���M�G��yG ��4Y���Y:� l��T��)9,p���x�eݳd	�\Yn���͵i?w����1��������Q�|C:9��|"x�Rا	,�Ǳ�',T�	�׳a	`JN
+��4}��.��z0v6 ��� ����Z[_&�H��ɱH�5���SQr�AV���a6��4��5���;��wH�[by�Aٻ��e��LA��_�`c�`߷PފK	��[a�,�>�Uib� ���-XĤ
$�6* ̣M��/X��*�T
kO)j�4���jklNs���U�`󇣨y�Nd�H(�o��,Iؑeq��
 ��aGu� F=l3����^z)��u�]�dO�S�Dx������ ��^�L��^a
d�Cy�+�c/L�+;6k$ϳm��ŋ_0k֬u�i�E8�޺��LO�TrrG $�����9���7��-F	<��p]�Qd��4 I�![@w������h?�F\5�s` �k��H�P�����w�R0:���^��Y�G)J���ݽ�b1?�r�dU��[hŊ��֭.ّ*�.Ǔqf�G~�=a
��.��ϻ�`���X�B��̪ �U��g�@F(��} �K�g�jx	(@X��更����a�ʻXD�ʤ�S`�!>���Ѻ��ɶS4���>�S�}G�1� �xJQ]�pRf-��DK�UWײ��Na[���i�O~�LĂ�q�㫯��������9s氜�裏���!���?�C��ȓ�2������%��ʲ;������������>C���D~�hѢ���-grOo3a�0nn��It���M��x�Lx2���3B �� %F�5��7��'d��p�@�R��5���������>%Oh ��K"��@��������˒D�;�V��$iܞ�����s3E#u����􉏟O7C��%G�)4g�?�|�(���������Je�ʻ�T�	�re#�j�GH�~N8D++�`�>ɏK���m�4��0�a` @�[��6/ۊ���Nx������G"�륆Z�/�O��9��V�����^j�HS<aP4�@N��>S��z1��� ���G�!|o���1c��y���/2�A������П����7�̒����@`
��P�ꃄ�M�I$P�_�XX|Z�C� ���{�e�����"���-Z��� N��z/>L8��s �O��#�|�?|c�#��9�0ȊC p�]5*��[��Q놁q�:�(:묳x1��s��N6�mI�%+\p.v�����7�N�����:=����F�l�̙{�n���xo�^}i}�c��4���(�d�s��t���e�roO�L�����!�����E.����Y�pL�9����|W�����;����;��Z3��E�E���g>��O���sB�P�+_�_���DnE�]�x>�|ұd��J�ko��g�}�&�=�jFS*aR4VO�
R��sv�0������a	�����?�����3����d�©��������'^ G`ta`
�駟�~l
&,a�����*�u���E��p�������.���-J) �p�*
��˖�	E<"v-��1��<���]�7��Q�b�|������x���l�=�k.�M��\0�O<��xE/��B�
]u�Ulp_���������׼�y�vut��W�ڶ�@sN=�.��T��W^�Dg�u)�kMYu���r��� M����^-�(�����s�����Lh���\c _�/k �K��cy�r�+.3���}5�c8���� {����L��,l 8�;���;n%�레�K�z!���㑏����7�u��]���i��#(��)��D5{^�}*�YL��3 m���C��R�8�́�b��~.�
�|��\�8F�_    IDAT,��<��.B�d����?:�.A�����cG�O�m۾kѢE_�(O9w����kni��T��g1���/Pm]�|������Bb�͊sM �����(�P�d���=v^�f}�H�y晬A��/}�G(� c��C�\�&�r$װ��E�o:�����詧�JӦ��o|s�3~z�����ͣT���	?�
�W`���79����Qc������k�>��+K9V��a@v�eÅk��8�xa}1�3�%E��tr�i9@8��JU�-^|}��'RWw;-�j=���4z��w��4}�!�(Faf重b"�%�����u���>��>�Cd�������±���+H��ԧ�3H�
 �z����(�ɕ�<�(.�!�\lf��������g�毮����}ϙ?s��ͷEz�L�i~�F���g�m�z��'�̎�_q�nZ�P���#`D��3k�,�X 3�%�~�1��7�J��r
_���cP���Q�!1J�%�a3?8���*<iX�����+_Fo��53i�U���L�Wm���9�M 8J
��(F���~���AKB�B .��#����9����b��$1��Co)=����	0�Y��~��[(�襆FE�_�Y:�#�Gt��W�SO�Ұa{З._D�L��'�1���Xq���L;���J���z��N:�N:�L��K/�Dw�qmذ�/^̑7�x#/�8�/q��%��AV=��2�H_��@��������~0H��tJVṑ����._1��ɓ�Ʀy�#&ͻx������${�q�]e��	��=�^~�Ez��g	���� ¸A	'��1�'`(h7�
��2�
`��a��g�i����aA�q<>ñ-Z��� �qMLAp���>�������t啋�����A�^��&Mއ�{�u��GϦD2Fi7J�YEdD��9gp��q!���Ǿ�,  �曯����	�vwSuU�/9�N��<K����7��'��iͿ�2�c�=��7ͬ��N��㽝��C�����А�v/^������s��	'��}��?�}���e���׿��H��={�l:��=��;^� 	Y���υ܀������G�����M]��
Ѝؑ_/Z���Lx�s/�6r�[�ե�3"xISt�!G�	'|�{��f�2]dK�%��������L��w=='�PBBB "Hii�@��҂!�8���w����f�$� ���)�؝QQ�+�9m������OǓĐ'�u�u��������_�~����?DfI'Wp.L�����Z���p�҆��68���"|���P��r̄�6\�n����^��]{�n���q�����[�ՕU��R/��1��� L����,C}��%�9�t�}�*�rjk-k��߫/:5�y��g5��V�Ԫ[n�Co=��`�V��4�<M%��7��d�~����[�DE��6��;묳�S�����'�ֹ�q��8�Xm�|7������8�b�s-�n��N}���3�ל�r7o
�S�V+�T��;�ν���L�8���=fӚ�z:�F.: |��O�y�[?��g�a��s��7AB��:�!�r!�)��@]��Þ�|�K_
�{��;<��0e p^N'�fr8�c�%�s1~�bHV��ٮ�������Z��I����ڔϕ�nMY�w�r���%Ӥ �f�$O~G�?�����k[�e+���^j�&}����E���Ƥr��^zq�~�����7M��_?��_���l0fHS���A�!l��	����)G�ڈ#�y�����?�A0G��7q�y���d			"�t YH#�P���+w�h�r79`���4L��JWM�SO�}�]7�r�)�WE��o9j�����Ӽu�1�1�2�������^�Z*�IPI� ��TX;�� k5�5�����Yp�q@�^y��9���<,+戾��t�؎5��Љ1�=!$-�}�7YU�	�Sz�!l	�U���P�{�K��1�C��ɪTM)�	��4y�t5n���!~m��P��FᕫW�Ա�CMMe�}��5mƹJ���Jjn��[Kڴ9�|>�Lj��R�{�q���tD/%���1�Ad�=��}�X�17`�%�!�c��v�i�q���6��"�O�+����X�ҥ�}>8���Y�|ꩧ�y�ۄ��L���wr��Q��lZ����?��,"	^�a���ks�F}���U[#��W�X\p�/�a�e�sh �EP� :��dђt�+B�q�� 1��s���}��� �j�☳(�����\k���y��[3*��)��kX�H�������ھ����&>��*T�԰W	����vH�	0��s���@�ZHh̨V]u��z׻NR6[V:ԆH�\kTwgM�T����*�Jg*a�Ѱyp*�+~��<�i��aj�[�xm9A�7���G bS�N 68;�u�ĉ/���f�,0	��h�+�=�F�tWOwg2٧�y���0~Ӗ�����yՂ���I�#�Lވ��:u�8t����3*vcG��h,����߀'�^<������9��H?�&��q�{�F�5? 3�����/� ��a���X�`SvP��s�)�8kz��O�k���BO��P�2���k�(E�rج$N��K.�l��UO���x���P;C�/��C=��m�n7ftV�U��[�m�*U���ǝ�7��r� ���BoAz�I�,[�kD0�K���#����B�0���ի��;��N���I<'	Q����w`��8��`����ӟ�e���V�@��s�D�Z%c�s�����xío�i���|׉�d-I-��d���Stҩ'襥��r�������z��:i2:	���Fh/����C��6`�>���SO���]�Vs��	6c��m|7(�F��6M&�N���gU��:gRd�P!��>U�V�V�as�ƍW6C�r�@�Ƽ��kH�%+i���Tʥ�%ns�fʪVzTKBrjjl����Xe�#U-g��ܤ���`��ը�V�K�
[454(�ӼP 8�$���2�!V�����,=a�u�5��H����P�j,�v���k+v�&Rۃ�@���.����j�J)˯͙3gp����_^�pT�<�;ߝhmjU�3�7����2���5��g�5k��ES�ދ 錗f� "��I�-i��	=���3_(ڇf��@TT"`��k,���7�d ��q�۵t�":+��m-( )_`Ś��F���QBS���QGMP:�[����~!�PS�Z1�KOH�FU�Ez�N������6��Qo����ViPKK�����j���z�p>` ;��9	V�z��a��s��F[�3�ӎ�]̙�� v��6mڴ�z&��2�{�F6��ɢ�j���}Y�qސ�k�H���ܹs?4�E��ћ6,l��6)�I&��/Sa��u�X������MZ�|e�`�m:�"�N�0��d�j��x�t1�`r�Y�pZ{?h6�f�-溸� �����v����^\[��|O=�;Ö0�P*�6B�Wo��a[���
A���Pt�^����$`^�v�>���T쪅H���4jX�O�Jgq�Q$�Qg��B�:�ڢR� %;��)U*�@��G# ��w0�����vK�-���~�^"�LxhBÆ�]w��#��v];��@���8���xa���MM ��G[Q�"HP @�v���Lx�A���ͫ4to?���A����2h��*��:�Lw�[C��@��8:�Tm^���/t��? ��cE=���P%��% ��DG`~`9�&ta��"��7�!8�=x��xƌ5�(�R&�m���eU,oWKKB�JR�}~�>��g�eK�������Sg��!~���P�Q�+����ROU�nӬ+/�9�P�,�*�H�FU����u�R���������p?Ha_(>0Z�����?���%�)�6u�z�Hڊx^�s/g�b����Ŧ��z�OT��8�_	_m��QZ�M�6q�������	£6�Z�Z�91�N$�@��F1���+ۘљg���?!�V� 1�s99k�g9�ҀNq&�t �������\G�������;��@��a�$k��w0�2ib
z�ڵe�
e(�פ�/n��ݤ��ʵ�  L���(C�A��C���%�	c��֥�6��;ޫ����/D���`utI��P�I�r���l�`Xg�;|*.��5~3���RO|3���0��~z��:m��!8�� ��?f��W↹ ��~��6 �	��b� ��x�z�Q@�����Y�R�>��J�mI�=eU�5�(W�Ѱ�vM�0Qd�'L� G~��� a�t����g{@�(qu&�
"h�9;��N:�t���(�	;N8~}�a�U*t���򸎞p�N<����Vuu�fUQ^p�*�*ײ�
E|�N�g̑m7��=V5pI� �b��������'t睳t�{NUcSJ=���,ڬ<�k�t�jh�Z5�T�1D �{��f�@�d�x�3�Y5ϛ7/�%����e25�1U0�!|��<G? �|G�	��s8߬����^�S$������O?z��7 VΟ�H�Ά����	�E�a(��÷�'���cJ��@g)��vT#XG8�e1�D@�|�^�z�i�:���	�Q�o�p젣��|�>��U�nҥSߩ�o�'w,]�U�\t��y�8U��as�	1�}4Ǉn��K� �d�KZ��Q���WB��E�X�����O=�mۓ��#Җ��f%�ٰ�'�!2��'���C�U<d�3w�4���js]	���fe������������q�iq���^�Y���+l�؀c�2�5��+�L��a����$%��b���d��锺J��nKSk�xd�@�`��~m����(��L�^��pq�����ý\�Ӷ�s�m���r;8F�U��z���ߵj9�[>�����o~���8L�����qoђ%�4����;�r�A5���h��{A�%�s�9^5oH���r�r-|l�r���f�ϸ��@���������G��YW�_o}�۔���Ɔa�r�y
q�3�	c�c ���A�^ۡ�����&�l�^��`K���ڮ��u|/�
�����*��s eL|o_�K#ĵ���e��|�I�jI�M��娘��R��j�.0�t��i�5���BZ�YPt֬�5�^�g;��m֖|g��� 3���`Ψ	�^-���S�W�Я�S5������'u��oՒ�k4y�U*{A�-ﳚ:�
u�ذ�V�N���e�탩>t��Ua�'L�Rʫ����o��)S���C�S����>����;5~�DQ��'_P6S�=&���B&,)��e0����j�ؗ?���x�k 2��:'�6f��zTŰ��ͦN������Lc&<w�����>$klX�c�$!jDG�Sź�y�j-w6��^P���ef�d�8Y�%����~I�Ҡ]�j5d�}|��ziɯuđc�����z�����+4c�u���ܮD�[��2�2����U�wr(cn_�ܡ{�	$����+ֿ�+���pJK����Y���i��>��Y�>������}�k?Ѩ�o�-~��;A������j� L6m}g�N�c����v�κ��{�|?��jb��cL�ܸM�f���͛w��g�mX�������
q��Aة�����}9�x��������{�Ś�O��������#ںu�f�:O7�0]�����3oԶ��pk�'LL�)�4~JgJa�!ޗow���^{��Y�A}D=]���V�w�O�M?O�B�~������K�])}�c���'ջ�H�B9��-��Y�9
�p�R�o� ��c9D�^��b��A�D�7�HV�fD������AQ;�ڏ�i�5ZK='����� �j�7��� �|�����UԦ�ل���ZY��=���}DUg�}�F�N���G+��t�����=�a�Tk)M�	O�4U����ne��yod0t���0^�|��?����jn���s�Ռ+�W�ԣj%�_ܨ_�b�Ǝ;A#F�JYJ�YU�4S`��r=.��)vְ����4����d���w�}�*w�-o��养ao�=� K�}l+��聾�0Q�'_X���_�����8�Q�G��jQ��ujj��UW\�amݒ	?�Z˾]���
5��-1�;T��OC��Ax��5Z������̪���1W.v��+��ھ���N��ܤ(�re�)�lP�R
;k�����p���S��?N�ʌ�k����o@�}��ڊ�	'2G$E��]Oe�A��(	��q����c���	B����T�յQ���RIjWt���]/<�^s�}Z�0�j�b b@�>�O��q��Z��S!�|H{(�Ϣ����Z�i��.��.�{�ijlH�ɫU2l���SU���^�;���K�P}#�L�Qq��6�U�>X <w���M&�;��S؄w&q@�^�r\_m�?8�b�����*�B�����+�iR:9J��Sc�p�j�&߽�iS��رG���C�O�@=m9�UkW�GV��!ky0�Imm%TV��h�v54���o?M�����&�"��ެ�z</!a����Ef�3G`t�6�[����&��:l_
�6�P��������c����'�DU�D2�B��5�kUw�08�F�*I��Y��H�bHN���X/6=d�ؗox���V�����];b��Ez��G�(ה�+9�J��	Gf\*Ѣ���&s�Z�[U��C"V!_	)�6E���PwQ�cn_DZ�c��L&��3g�����}Q{y���RQ�QwL����C<���ŀ��.��xa�I9lj��m�`�d�lZ_�(4Q��0��,���5hh�	Ke%�)M�6Kcǎ|� \���9b_�١{�{	�/[]�rc��Z���
ʦ��64��O�y�pr�a�XcsV�JU�JZ�dF���1~86�ٲ�������5@��s�̹aPA�^Em��ƞ�I�L2�L��</�&5TC� �ɐ�P��o�+�;x�I!s�d��x@~;��Kg�8l�b����f�~�xPU��������[�D8K��̏�C[7n���w����jZ�jc�u�$`U��-;c�<����b�	�\{���^�������*��C�Ր��!#JE�4�T-ըc�9Aox�[�/���w���Q�=��!i�#�N��3ژ�$V�)��u���%��9B��;l�����z�	�wY��Xs�1���Y�={��&MZ�'�m��	7���Q��>z@�vR�Г`��T�j�j��/�Ԙm
v(�BH��3��������s���:Β3�v�˲c����]?���7[-M�ri_���/&�eIԣ��uИѪ�s!d-�j�ꕝ��;U.7���3�1���)��פq�C�{2��ݟ$�w ���Z��Q%*y�SE���t�{�PKK*�(���`޺5����a'�R1���ȐmZS1wg�1��/~1��Lc�5���ט��Ǽ�{�����=�'��=�s^9������9(F��l^op  ��ٳg�8� <fÆ��ʹI�b.TQ��O�TT��U0ឞ|p�F��|�^.!I�����`r�9��zI��d��C���Y�X��ls���F]uլ���	����Z�ڇ�4rTZ��F�#_]Z����}D[�$U�5�k��ڛ�\��1�����O%�`fL��l�j�_����˦{t���5u��*;B��D�U�JV��m�-*����ԔN�����ZNJ��u�� ���BJR�<x�8��} n���w�뚓K�� �WٜK�`�Sٍ�c �[:ǳ�cP�R��R��x��M�8��=y�d��|����S�7M�6�m8Ԏ�]Y���*�dGӱ��%U��=q���t�P*�S�3f��k    IDAT�6iX�,y���Ջ\���Z���g͚����3`�����n��'���I��q�^wp��wvj�҂.��fuw��Zk
*�	��P:��VJ[ޓ7t��	�q�=�ϪV:�ؘ׽snԥ��T2Q��=�\������c4|䡡VwSӨ����H��|�+�O�	�1��l�%m����:+lr>XCUF���!���� (�&x.�p�����JYj��fJ��ZĤ_���a�fV�v�̘�+�J%�L>����4� <f���M��IM쬑/&�А���V5�4��'��N� �@~��0A�ri��v �E�@�)=���?��E,%8�=,���6wxGf3c�-���؛8b�QJ)ו�,{��t��g��NVk�0-[ܩ�fݦM��� \�ԩ�â�y�:d���+C��	�W�Y���>��6���{�����V�����>���UwwR���7:�ȉ�犪���S2I�r J`U��Ļ�Pj���
PdU�R��}�[21������� �ls��U`|�ƦL�(\�l����2����N�j�
?y����t��n�Y�	{�mG�oZ3���cgQʒ퍊ł�M�)��]��rZ�	S�޻�� W;�EP|:�DA�z�O>�d d�f��jh��m2�T��v���W^yE=@<�x��� kI�[���KK���Ԣ���7:���Ӣ�o��iׅz�;@xGQ�T�h�8�����K:wH���K�X�D�y���m5"������s�Yڶe���S����ZZ�wާ716�0cd��u�H�����  l����/�2�l�.��5��~0�x ��am�q~���N��g� �"�`��^���f�@�� ��`���7���~����^�ʃ>��Ae��m��7�t�H(IC�I��]��&�]�>G�-[��q�lH��C`T8�cMf�(l�6�c��^����4/�v�P��P��[��V�F���"Dvr�:ur�vI�`}fI�ۺ4w��Z��Eez������3V[�t��SU(4�"�	�{�	_��L8קþώo���=q���?J`o
��¼]0�a�6iԨ�n��Z]p��ܾ]w�u���!�����Ə���C��r����|T�/�~������3���g�s�'?�I��:ʁ�������^q-r�6N9��ٟ�Y���e˖ ���`��s��ζiv�`�
̨�<�LX�C�= �H$���'>q�����7to ��ܦbG^�v�ο��=f�^��"�Z����P2�A(�Lh�p1`�!��ݖ���ǵл���`� ��t����p����aՠe{CM6�+��<��CT�@ǖ-���}J���Ot��-z��������/,ѕ�nPG7 gBhM��p/��,�K����N�?E���m��u����Z�r�.�B ᖖ�f���f̸@=]ݺ�������:\7}�M:�4u�t+�a�	".=����6�\����
@���؟P@�`[2�U�\o�����??`&-�9:�@�U�#��3��6p�o~���S/�+'��'|��[���8?�u㉙lJM�-*l���<C���4����Z�z�:;��	@"0���y{Z�����#
+��1� .����f�N�%aI��,0i>f�ZL3g���,�ӯZP��Mw�}�zz6h����ʫ.R���z�՚:�usD�pR�DF��my�8%SDGTT��ل�h���x�D䭵c�ks;gm�w*�\d;6�Hj�kCk+W���gU
ݡ��=��W��|���o���-�'���l��#�Go�t���J�e��2��0vWp��N~��O"Q�!e�(+p
��7�b���WVӧ�v�N>��p� dmN�M�.���:̥�.~�r��`�t0�(���N��<o޼[�&<b������]ԝ�.�l�|���/~���\�� ��h��.�(<���Tl@����~W��կ�0m.0pp/<�쪊M����Z�e�8�aq��;k8��w^�d���o_�!�������MU�	�\֡)�?���&U�TQK�p�@��{��a�)6�;J��1�����"�����|ò��=��(�L�1�Z�?I� �l�r=���Ky��U���/{�e)QYL�w/lҢ7�u��S۰����Cj��ke%��Q'P�	������}V˄��{K��r=�~�<s�k��N�0hB�p�a�4�3�5p��
��/|�g�������o;���
sD*���}��w렂0!jlX�`��'�+EU�5�~̡�����m���_�,DX�,&L��g�5�uv	�H�8r��^�9���P}��![&	���/gZ��bc|l�Ahl���}��f�;c����9"��L����ש��M+�nׅB�E55�L�P;3J*�[O�7����ncfj�J;�vV����WVT|�跗S�����u�ܟ&�P[^��KC5�	ko��=KS���&Xn�r�mڶ������{�3�bK�L��(/W��W׀����0����-�?�;wn����W�vj'� e~c&��=���e�L�6-��f��0�AI���9��7�������L��G[X�s'�Kj�Z9�J}y�A�����ױ��-�Z��;Q3g^��|�b�k�7�~����+* ᥮�6tA�����da�x>R;� ��.�(�{�����6D� 8K^ ,!��$��}�{Ò;���	R�J�Q6-�z��mXV�|I+�n��om��S/e��׉�6u�ƍ=��9� ؄�|�q��+L7���)F�x����7d��p:�$���;���>]��i?���I�$$kZ�j�>:_���F���_���91���
#�+�ʹG�\���L�;bya���as&,��/�g��v�K.�$��(�M��ډ'���ް�x�A� T�;�j�S܇U;�8�29�����=�d�9�;_��v}f���D� |��'��ߣ��ڼu�J�r�	�����j�%9N?��p��A�'M�:Jx�w8����s��9�ӷC3���p�eP��=�RHX>x�/���� ����3�UWG��Ŝ��)<]P*1LK��UCK[HJ񌡨�� �
	��W˄��m6�2���"!N��>�]6Vf�S���
����r�I�^d����	>Ԗ�_�k���{X�BV�ZE�N����o�ӓ+��Cޠ�O����R��U�Pϐ��V�Ř����g�������k � I�*��m�g>��w��L�iچ)@uL���� m̞�1��8D$q˽��1��=��s۠�-�^��ݖ)����E]�����Z�zE0G ¼�����$��!cǍ3T��a�,3(t����2�����-\^�C����͂����aN�EQ/��H���PH$��A�Q�@TG�
�j��ɢ*�h�:Τ��I4�^��L�]~����'���z�:Q%����8+XA`
r.���1+����P�'	�A��%+^�#_���ڕĴPٮD�:UjUe����:b�jic�܆����)��T��ѕӜ��(+��0q�_}��!B��9��SO� �c�k��� p�;S�8c"�i�c��ۨ��<�Wp����q��3��
�ͪ�w��={�-�
�0�Q�V-l�&aFx?J�_>C�-��~���X��P@x�ĉ !a�Ȅ4�S��8?��9����`� ���Z�[Y#P/�]t�!qQq�Hl�@�uf\Q�RԢſז���I���H
xHM�����J� \Ӕ�3��Ã �������~����]B�V>V4f��ӡ�(7!���q��4����ڐ�Axպ���IU�傚�j��u'X�Y�L�&L���*���9�&\VR�>s ����ς��9⪫�
�"A�0����>�g�� <s\�0O=���Kd[3`��ò��y�
@�{::\���b�zI�O�}�݃�#7�\0J���{:��ԪCF����J��.���.؄q��@v��4��q{����YN����l%�&�%�� Ll<�=�%��
�հ���̆�X�����|n�~����ٱ-���
��4;,zi�jlł�!U7GL���^N+E��^�1'-O��񋱩Þ\;�,[�}���^ �d���V�3^S����l�X�f�}d��]R[S�ڇ�Ԑ�&��Ҫ�����>H�}�:�����@��WQ��	��:v��7懛o�9���8��l�Lw����50���
��|�+�r�����(!�S��p9n;4�`�&�����L�"�&�V�~�{�yP�	S�}����O���H�5F��ݺ��[B����%55�v��O%��a�6Nl,��=��H������;��܀V�		AЀ5�<0;��0d�H�6Q~c�L���jG�T
�Aw�>���*�rJe�J%�ܯW�{�B��I�T�M��d�: �y�;�#����8j3[�G3#?�o���f�^p�|lj�o��6d�(0;��"��0#��]���-�J���%����0bs�����Ǳ؁h��a�~|��!�����'c�o�e�p��WHV�nw�3���{�zEc�eD[�N$`~���s8�=��8}�m�A8��Ǟ�O�?/�}̠�7���dM+V���?�\G�=x����<]|񟅚�L�
��R�vmڜS��c�=��R�=�ݳì�L�����7����I�/D"Z��<���{�a���+��2� �I���	�x���L���yLÜ�aA8�o,��p:�~��{��Ƞ�1��Ft�_���v2���������N:F���i�˛T��sw�iϧ�;�&�'8��d b�AS�>Oh���_l�a �����*)q4��>8�x�Ax�ῨJu�F�H�o8D6����Y%z�5e�5�盂3���$l�퍨'����%�`�������	I�\�;u9xI'��~����'��<ϓ؃� ��������!;?׬����:l��\e�fE�wo�j��~��ab��z��������4էhl#7�������0�8��Jn�{B�
.vj���2�ǲ1X��v�ڔ��ξ��&������^���g��n��ݯ�]�A8����ݥ�l�M7O�ԩTQc�5dҊU�U(��N��(-u�&����=F�.�>�\sM`�8�*�[�2�����o�'Vӄ��^����&�6K �=��9��Y�C���>�{s�p*��ڽ��{Ӡ��ȭ�6�t���ܐ��O��:����i�Q�!��~�֯����^BG~tfANU�0�J�޿���&����� �����n#�'��3��L?!z ��z����|�T��%U��o���ƌi�{.<C�-���V,�Ԍ�7��3�J�Y� �鐬1n�X�ӕ`SN�2�k�>sG/H8���qW}�9^5�@h6䕀��`&�I�Ak��{�fñ��@36+<4?�7@���i{2h�1ӴYē�>���ǌ���d�x�?Ã����m��=��$���f� �^_���&O|'�� �qj��L�tr?ڱ���឴��oF��gE�1l`������"�?׫�6� �Y2�e+Vh��_P>ץ���u��v��J%kھ�����J=��M8���%�J7dU,u�S�EdU}{4�.ή�����#��E88
���г����c.��� �ؓ�+�>���w��x����&L;�+˲w�� �9s�|h�A�mÊ����I�R>�Ne'�	�x��B�U+VkѢ�B�bVeA����d<� )��x;��^f�)��{�qR�@h3#�|�|�p���\G��N�Ɋ��-�}�Mںm�.��}�P*����AS'_�Rq��զ�-'�5u��^.�F��pn%l�֎R@�xbz¡L�rI��X�<�e�cv��;E܊�l��f�?�gGGxBs-��خ��������0:�ȸ�eO ���cFƳc`5�5Hr//�<.��v���\�UV�0��0�Y&6�+��9�g3٘�ǀ��C�����y�N(B&1��qR�MQVj;Sd|O]��c��(�X	����7�Y+���.ї��E康����;��5����ݟ�>����6���;u�o�鰠.W�\K)Q��Q��`�a�q�	s����� D�^�+p��j�z�������I#��3���๏A�d�c��ް���|�+�1�|Md��j �{�w�AxĖ�G�J'���)jGx����z���j��	ڴiK��X�[��n�@a��	@�{l+[3{�mz�'OA��9္1Q<�< "�)N=��}���i��c�|�����sp���?������߭�{�3K��U����9������ՠ�U��kRO@�(^@�l�p�h�P�|>������sO��0P<)~����;6�&���`�b��1�`�2-	�=/���6��|h�%��Y%�4�q�������+f�1��;���.blvn6�d�-�U�Q۞m���� ����l�1�s�e+�X�Ǭ�J�כ��m{��?~���to�0�{i�b=����J�iB�c�.��L�x�+}����<\��>W�&�j-�r%/��Jg�D��)��i;~�O}�S�= {�>x@������n<_p�"#c��Am��q�U�My�����}�k}�����d20��	صaarۦ��!j՞��U����9g�+쬁p0�tҚ� ��a9F� F���G��أ� ��3L�a ��uυ��	�e��}ܽS&�H�Еל{n����<8�?q�N9��\�E�ϸ^]]��R�0�z����`U��8ᘭ�^�!����><�]��s��ؽ�I΋Ɔk扣�`�g![��#�0}˃ev��1��ywț��0 t*Ê�u=|-�=<�hǸ'�N��`r�ެrP4g<�Q{�N�dblfMi��oȄ���p<�|�mA���@l;d��o��(װra;|	y1��o@�,�y�6u��ܗ��/m�r���ݦ]�*l��6���KȌ�D_9��pQr���h�s���^5�AZ�)�	/]�D_y��ڼq�:�A��1K_r��nަ믿M�^ت<R��:��	jjlS��W-ݣb1��T�T�;�c�W���r3�3�hcҀ���`EO�\ܝ��=8�Y!#gV|�Ƶ�
�W�}������J�8��MSƠ}�8��6MjimJ��A=�l6�|�G�R^��mz�����x>�T��0����[�D��v
�U0�04��ٌ�k�[x+^��`�;�J����V-Z�s��-#���V�;�`-]�AS�_��δ*U��l�Y�t%d�%zkg�� ��b��&K&�MۘD '��53a\����X�Vf"�6@@��&#�8�}l�o�c�e@��� �k1<���J�����asO�E��,y�|��2�20�7?���L��9^�܋PĘ���'�0�xc��!��u��3q�iE;��ל�In`c�"s+2���Y�Z�f�~�����O����˸�Lm�9!� x  &;r����f���`O�#<�c��2`�{�����{�a��J�+���/�1mݼY�����g���g���C�7��S��TÆ�;�Oo{L�W�T�+�P�,YI�o�p��#���{�+f�?Bvf�V&��.�@lvd��EE5�-�I(`wG��G3o�s3�W��
3����aЙ0�a����*I�9loT��U͔�ΦT.��\*�
��&f��P��섁��!����N,x��`�R�����6U�.>3���F3�@��9o1ס��Y��˺⪋5��B��U��1�P��ZkP��P�rf�m9�
gP�>�cS/����D����xU1���ٖeM��FN0 �6@��D�0�,E �AD�p�m�n��&�FG���w�sv�= 	���� ���$���0(�e��;�0��m����?rR    IDAT� �.5�$@6�H�#�8����D��y�| 2���(@�〓MA�=��g,�8�������_d�,Q���x��w�Mڏ�b����}u�
�!}8��2Gބf��b��ܠD+�FI ��I3n�r��(e���嘕;�2xG�p1���|}��|ɲ���Ǿ������G?6C�/;7���������Rg������c���X�E�=�JT����:���y睁�!8"���0����u�Y�>�!3�nPzȜ1땵��e�x���/��(���J���;w��wܚ=��.�7"Dm�5ZK=')QM��= L	�r�j*��s��t���C�����W���IOL�����}�{�+
�Qs}MlɽA�>���x���0�W����t�k�J�lo���.�x�&L�d��&�t2!�=~�{�K��#a�01� L@��pfr1i�����a�ʀ�=��P���z@���I���	���c�� l6��� Y �s̑h���1 �`E�\�5v(a@�~�=?����o�&�p��$�� 5�gs��0`À KD����r$%� ��XI�=�N����
��K{9ӌ��� "
�����;mQ�\K���w��><��slR���{������	#o���j�%��! >���ڦ������ %B�b��W�����0��	�^�F=�9U��P��;��%�OWc6
�,}iS����o9N��c�N��L֓z�+��z�I �E��<�9�E���>��I�.�߻����~;�/$��܏�?��>�����tz���8�L������}�'+QM�)��� ��Hk3/�c��߱���	 <ӶI����&<Px�[��%)٥C�t������s�\�~��m*�S�8Κt�%S�Ru��;�^F�O�τ��g�2alo�\��Ť�@���yLT&�w ,��e��4|�? �hh� �0T 9�,�̓���n���И��;u}W��r��Afk<&L;�:�-}x +,f<@啓��PZV�6#01Q��s�o�t9x@(7�%���\�yȁ������� ������hh��=q3}����N����ʂsQ��$����F�|�c���W�[���{�3s���y���<�N��������Z�2��� "]�s�ua5�ɒ�ߣ��1��Z�f��ŴZ�G���$��)�TO�g�#Ko��1�)+��aj����x�m������[1 ��}����������9��`mM����- ��=��5�����@U�*=��ڤ�LM-�xZ7��Ѻ�=��޿UWGU�23�P�d��u���J&�}��uڶ�6j�E��<�}g�0������1�cخ�� Y���f�_& ��x���ȅ{���]Lfl���
R��"��59�`E�����1{uH�'6���)}`"��@�z��cF�@?m�� �d�� ��}z�8����N
Ϡ��"`�N� ��?�����x��ov~�^0_�L O�0p���C� 6ރK�"G���PJ���D����w���|'�ŃLQ�(&@�U�G���x������A��B��Y�)�}r�(VS<F�����A��3�/_@�1�R��w�:�4���Q����˵�2�[�U��������>���t�Wʴ�Ǥ�v���-�ܰ"�jثgcW��A>^M�'�ƠD"��x���{��?�=}x�������7�o|yA[���;c��t=: ���K�8|� eM��������G{���L���e��FtC�ح���GZ�jE �r�#T�K&��Ғujn�\��i*ժ�L�,LB�t���m�"G��
/ �2��ق�2Y��a��b�9
 `��Ra;aW�B~LP��L@�8�Cl�+���x �XI�T /�`�8�X"�	@�vp-  �rm��.�o�\ c p�]�`6�➀�}(���>� O��p-��<�L
�8�@�D! s�N����(-��= |��ʓ�Se�/rfL�f�N}��<���Q<�����E?�/Ǒ?�@��q�, �ǽ�@�PĘE����ȇ{�V�y()�j��1���x�L8U��W�s=�J����4���?�!�)�F56��ط���y} a�aja��w�.#[V�����$=�-�=���������|��0�o����W �9b@�p̄-�X(ql�;��`�'��.�53��¬���M�Z����,VO��`#.�XK�VmU2ݢd�Q=łҙ������:z^^R�+�/��b"���y�g��� jdò�A�#��a1�3a�,���d�������^v�"����y�,���4��1�Ñ6�7� ��`Ұl��؃]� F&|O;x>��P"+'� Z��A>�>0=;!�5�{1�A��N��L������	
��<��� ��1�hE�;�g�F��=�����M ��G~8�������v:���
�˸�Ǭ���V,���&���7a���٫f©������W��^SK�Q���U5f����c����C_�lC����+W��)rʦ�;~���66��fKc��{��,����8a[q�����nG����>���'��<ۥc.b�;a�	;��>Y�(�X��,�=i�@�Q��9��5[l�B�U����K�
�'S�+�)6m�-J(�|�T���C� �ђ�/M���T���d��H��l��fb���m�LjX8���o�0N�Cc�����M�q�	� ���
L`'4�&�X�k���8 N� R�t����㏶�0a��&;���P�PnY�6Y�{� p�M�<��w���:~����y> �G�0\��=`�0x�J�N>��c<����L �D��6�˱�$ Y E�B�M��6�/���N�y������$��߀=�����3pl"_��&.�g�=9�ӤdwsowLx��EZ��/�g[U�[ڔ�^�D"��l���V+��c�S&۬D�ݐɈ�nM�R�~
�a��g�8<�]�a ��@H����ڑL&�}���_�'g��5Llnp�t��}a�@�N[� c��Db��B���*�.���׆�W.�`�-R�M�>�LI��
�dB	�K/��	&*��Q�x ��0&'툵:@����6:6�D�c@�L�
83��d� u{G0��� �mj�m��^  �( � m����Y���B��m��eN;`��
����W#V�<`�9,�9F���=����8���;# �6���,w�#'�8������w`�7� � �ڶh34���_�k@���1����]�lA�]L'� xw��w�8oLP����L�h2�{s���=a�ƴ�-�w�wC_ c��M�3C�v혫i��z�G��Y
~��ڪa�KJJ��J%[՝��w�Kc��J-��
�j,��|h?�/+{���x��Zy��Y��g��a_o"��&�zd�Θ�>��^^�Z��it 3aw¬�,ƃ��owfwygߛ}9 ���Rʒ6��h_��Ɔ���-jmI����ư���Et�-��'�T��Q�]M�K/	f�x�v��ba�LL �� ��9*�la4�0,�kP,�c��!�����9:"L��ɲ���.C����� �a��	 A����j�e�Ov�q-��y�U����jh&ǵ�����h�8�u���9�	���̑��> {�Vڂ����v����z�'�B��.�ȹ��YA 3'��S��>��!|���Uy�p�'�w��5��
�}��(+l���A{h�c����Q&N�F1V��`�׮���#��\�*QN*�����/һ�}�ʤ���%57�M[�U��A�0�*0ߔ*�Bؙ�J��V�N$���V��_&>�3G0c�F�h�O�7q���}ʉ�����M8�>�Z+'H[����D^�t"�	aa�6w��Zd��A,6Q�K	w>v8q��߶+٫
��5kV_��_D����R:��a*W�����M�^�Ӫ���K$5u��!YO0[��j$�ι�3 s�D9�1���Q0#'� 8N&�3z8Ppvru(��ISbr��F������@�k�T�}�г�Ӗw��A�w�o�D����>�
��(�X����l�ٽ��x2�o+����J7^aœ<fJÞ��<1��m�W��4��� ��noq���w'�px�ɔ/["�Ւ��N͞}�f�|w����0L�B�::ڴ���̳��z�I�럶ܿm�M�(J��Ϗ�W�摝�~_~W1�M\�E�<_8���=�ұ�7[��7	QTs����W
$k$ʥ��eBD�!c{h��D��~��,�����w�b���$/ `qzk��⥃Y@�]{�}!j��j%�[����[��z����Mo�|��߽�^׾�c��ȆR�,���:uZ��T7��?;���+�y�Xi��/��������7��A.�,��c�B^^��)�tt ���q�Iag�.�R/+�|1 �n����w�;c.���o+���p�T�190��0�K,�e߳���e�6�N�1���_�|��+�݁���k���/H�����{�L͸�\%Sm�Э��vc�KG�=Q�v���X.)��(A��2���!��7��x|���v�ج�I��q��oכ���c"bR�Xi�!?�Ǧ3f�i�`\I�Rߜ7o�5Nػ-7�;��\����p�݉������f� �M1S�Ϗ'M�<��3 ���ۖc���`iG=a�t&�c����G>r�
�����t��h��az��՚5����ި��)M�2]G�K(����5Vvd�ē�6�Y�Ď�ͼ�8�.vDY~��Ks�-2`I����Vlv*�go�Ҳ-��F�d�f�?{g@П���Z���u���?>޷�U�p�~�ցd�������$ f�Ⱥ�.fx�] x�X�N�>��s��Қ�w����g+�N�����>�����ܷ��}�4�t�
ee���)��L��vY;��äͲ�j���z0�8z��m�G^�7����Y�Wp�o�m'�Y3�2�4t�p�o9p��έ��)���90�r��R��J��'qƘm;4par�`��U�i8`�q')xpƬ!��v,��h:�~�q�мf̘�g�'E ��T*���>���~���М�7���&jŲM�r�z�[T���� l��[+m�i��;�ENQ�ض�	�d���,������5��<�cVX0 �M�K���1V�����+v������x�����{P���3���{�t���9�+6������;�>0��uv��l�*=�p��][�>��;f_�K.9C������}���i��7�;�ao�r��a�M*�����r)v\�v�j�oV���@إO�`��ybY1�#�1��<��.��0��8̔k�)1�ơ7op3���ǎ�qՂ�bω�0�R�+J4�B����`� \Xv�� `zY@�܎�t�[&���2O"��]����G���Y.��eĪ��y����Թ�C��{���(� ������g��eK7�]��T�֮j��n��}L�� �΀�ϵ�����x��) ��o�a����l�f��2�HM��g'�#C�K=��\|����"�������s�q�������̹�;���|cv�/e�kNh�������ڦ��U�5{�.��Lm޴I7}�.=��f�s�n��^�w�2#���Xަ�Ɣ�lWQ�9�CD��x��ؔ��31�`�6�`���'59���qm�o\ɐ��T���
ګ�}
��^wۑ�����jI�".������	�1w��G�XK@�Ѩ�P���Ll�r�=���6Qx��tU��Fx�/����ĽB���#x��Ȅ�ӧ�4:��:+��f�}���K1�@}�ԡ��ŋ�k��7����0*(�p�c.TQ�];�\n����M{y����P.��?Nրh`�
��7����6���r]7!vJ�m[C�.�3���.fb��eg�����
��;s,�a�1��@�1���،gv��0�=y�@�����X�Ǿ�@=�4|XBw�}��N=G۶l�'?��?O�B���ןt�&w�����.���T�ϟ�9��V�g�uV�%|��I:�EH�&���*~�6]��
���́6IX������+�x�o
��p��/��?�V:�P̉>�m!:"W�Vsk��1N�&�4������fR#DK.'.�j� ��kw`���s���XQH�#�"�ŕ��������xІ	V+�\���wݬ\n�.�r����^���j��k�+`nQ�<u��7^rPB������`��c>�D�����˯���8^�}�c}_~�
������]:ۋmZ��$��企�lo�lw���-�8raW�tO��33���	{��}q�.A8Y��K5�#*�t�m�t��4m��x<�̏�K���ϫXn�M�Cc�zk��L$ECM�|��ɺc��6�c����o㋽�\�H!| 4c�ӟ�t�W����^�r.�?ĥ�L?��+Lp
�φ(��'��g3o9�5M"&���y���e/�W
'����\S��.��l�1�Mԉo����B3)�1 �d�1��7��v!t��Ht�����������,x��~z��E(������}:ċ���{lی ��u�?����z���*��V�\֦E]p����;kXKk��+u�Q�ao!}�^Lxg`3[�#l�I��[���(�3��Td{q��7��F9:���!�A�n��b�pVK����_A8fJ���f�x��&�3>�M��?�Y�'����p�utDM�V.����/��-�[o�����U[K�:�KZ�l����s:f�)�d����^B�j!�Q�^g#�	�NoBxΛ7/�ѯ��}�帆﮾��0���6[G�x�ސ-I=בI�8Nn�w?����0�܀2��duȜ���w�sO�{ｃ[�}��|��Mk���r`#J���:n�&O�4�5��z�kO\:n��@3]w�F���R�� D��sx	`
�E{}�������*0�_��^�Č���5aK�n�uޑl�7(ky5d����!�Ӷ�5�6�Ce��/m��_�B�AU�Bմ��M�RG�=��~��� ���۫ /�̈��_�r1+f���Px1�s�u.C�����D�_��#ݛ��}![O|�W�Ǡ:��&3Ƹύ��Y2߹nn�t�K��I�q����jǽ����@���Ym��HT�l�-\���;�jx[Vw�y�&O~��U|ERcS�:��Z���9٘!�t&2n�[��l9JYƊͅ�0E�w�y�}B*,w�����׾D�P����c�g�F���1�l�u}�wl� �7���T~��D��H$�Ycp���Gm^;����6��ՊԚn�ȑ#t����[�<\���9mܸ9h :e��
B�|BM��}���q�&�Ɖ��6��\�i�L.l������~��9T���k=>����=��Y+(��Ѷ��LKɜ2e5-_�]���W�6��%K�ӧ\�qc�V:�Pg�$lP�g'!j�����p��
�ūgG1m{���I��]��w���cQ����������TzE�?�0fz1 ǡ��x��α�|g��ګ%?�J!Ί����
�^��db�;�=sĪ%z싏*�ա�mM�|��:��w(�%�?���(�fK�����$�4U�i��0G�2��~�0'xS Lv0YL 8�#�3\��?��`^��	�ZVvA�ۤy�vx��5ϣĀ�R��3�J}u�w[�GoY7�9���D�sò���t����굫�Ң%!D�F0�A9f�Ih1j`�y�駃��n�Pb���g�}v�� S�?�q_	ź)�\��2�X    IDAT@9m&Y`;4z�ZT�ܭ~�_�e��P��L�j%�Jy�֯�R2դr��Z���UM�2K���t2[<�w�;[�ƀ�h�]��}����U�d�oX���۹����-�����@pꩦ�o�ݫ�	�fY��������
�����n���1��Nc6(�~|3�o�
����_Z�HO>�
�|�H8��U�ښU�w���g�E��S4z��T����O��a�k�U��W��v>[a�'<�|�M�b �܀�9+�&H��"Q��b�\l�3�����e��C&|Q����:��>��~ �<\�����}���!j�L�=�#�V�P����r��k+`�%ځAb�o6��/ɻ1���л��J`u�%xY�J�_=N0�jQ�D i@��E�=�b�SJ��[TcC��96m	EH�	v��	�w����
���O���`��'
�=�<���v�>|G�aL^A��v�mF�Ն�ӫ�����A�w��]k��� ��x0���!�mG�kT�p�!ż��n��l���۱+Ξ�#��Z������խ�tF5̉Y�6�R�*j�*V:^�)�*I�%=�L@���U�Ʌ�K��o��P��F�]�>�7laFr��3�-k0�)l��X��vk��W1��躐�ìA(�O>
C�,V�U@��s�νip7�����#7���R�>&�9��чh֬+�S����j����`�A�F4ڱu| �l�6��BC�N��`8��s�	ڎplϘ%0e0�|� �y���A�~~�ew��\T������B��v%��'WS&�Q!׬tf��h��.�eM�
c��1s��s�*��Tcd�l{��cgVe��5��U1��펾��ڸ7���L�;���<ۀ3_��ݫ}��n,�X�Y9%66),��8����O ���Ήw�v��/b������x���{��0s+V걅_R��G�DM��6e3 k��ʨ��j�����<\�dJ�f���3&j�@n.gi�1��v�m_(|�s,��{�E�k E�E&&0�|�6��{G>�]��^��^�3��Z����o}K�j}�@8�zjޜ�T&Nx��� al�8�ƿy����*=����_P��ҫ��p�1`�DZ�P�`ԟ5X8;/��'��h;�'�k��&����%�k�n��>�9�X��oK�͋E�|x�9�C0�Z5�bn�~��h˖5��ra��d�I�|��.ݢ$�Oq�%s�97}�e7�(��^		u����&>>��g�"J;]��Yml汼͢ݦxij��g]�j�h�nWv���y��f�՞cZ��#O Z��Vef��x�j���6  Kq���{��7�
Kwf�**fz�{�$o-_�Z_����uu*�(���M5�;aӃb1����\�g5�ua���sy0}_Q�|�P�����sa�l.K�m��"?�l�!�L���k�{0�T�՜�1�����J��^�rh��v�S�$��ٱZͤ�_���9��[�='��|�	�8�m�2e�~�_?Һ���UQ��8�H��e;q"6	`�A���Ʉ��B������ H�~�,� �ܹs������߅R�/����c�?���h��$s:`L��s�C!�l��_آ�n{@[6W��XJUKV4m��z��`JKb	�e��}���~�~�V`\g���o�|�X=�|����	���N�ݱս��1�}�l+�x%�@�(��\��8��e��M6Sp�:�*���}ضH�0s[��"���2�\}϶a�Ǹ�� c�s�&�zD�����]�)�]�A=���/{g�wU���]g�Lv�UYٷV�E4 	���
QDY�E����Z�B
T�.�V�\�hA\ؗ���$$�}���~�?�p�w&�dk�:וk2��_�y�s��~���tw���m�矡Y'q�`?�g��Ʃ����^R=[��|~�����L2��eW9��,ކ�x#&]�5!��"���� ��c����
pSmyĆ�棵LL���B���;{��%#S�j��$��h4���}W\�ы�����;c�m�۬Yvg{��P�lX���	'�E<|�֭_�j�2��V�a�µ_�:K�P@��\�a���p Z,�����ٳ����a�qx�OX8B(�]���ج��~��5( RR����T�s��պ�y�K��~����������k�<�0 <C�75����k̪���1b3d����1���f�1���m�ɏ���A؆(��l�l�F�G�4p,��F&8%Ly��d� Ą�p�Q�b`Hb�f��6��*� |��q�et���@��������>�a�8��%r�a{fɳ���w�&�e����B��z���n囊�h�:�2Z��/�`�U���Ԩ'��S��L�a�q_�Q�>餓��#E��z�	c+�Py;��
�L��0(�
��, ���W�}�,a�p��kO`��+W=��Q#&|͂�;찱;ވ>۬}a��Ca���3�x�	����*0a�#PBvj�v�Q"��'��}��G��k_��`�m������ �2�����;/�7HUÅ3���s/ ���q�W(���{nծ����9G�e\����^X%�z�T)OR����蜹��mӶ�1��%~5]�6�R3��و��04oAgl1�\��צB�N(�3��C�(��PF���CHG2�i���|�.�B� @�>3�a�� `�=6�iO�@��a#������
8����=ٸ�~���"��T^0�]s-[Ӳ��ۿ�j�&�gt��wi�i'h\���ݫ�>�L?��ot�NҤ�;)6����2�����Q~ I��:�������pe
HiE�+Ű���½������� n�̡d�_�	��˹�������g�;��5�S��V�\��]{��c^�rʺ�'�ˇQ;�z��춗�<�=��
����z�,�a�q-����\�b(
�b/`�-���=��&fl��k�b�$V�1(9+�>�Ɩ9v�`u�����2����e�]�re��~���я�7��=ۥYo;G��dU9�)+�9s� ᰅ.)쾙y�[���� oW�3kq��<q7�.�38b*.�v�7��"
rT<�_���/ڋ~9�;�}f���"�O� ?���7���'��nﲱ��6h�͌��f��\����������s��v@V\����3?��Q}��E�'�/�×�Ws�Y�J�~���u�u�V&;U�/�V�L�_Ŧ�����BzA�L�~D[b���7�����v�ϥ���'�0ǹ����d��0@�X�zꩃ�`�Ƚ�,��(e26�F2*�q�\�*����Ύ�Ps���c
�u��v��q��ÓڟE��v�駩yBQ���*��I#Q���q1�:��RlmF �hX�?��?�O~�q��!�j!t�q��^��,qA��dל'��]c�� �(uU�L^=�}��k��C?��{�����N;３��J��K��UTU�h� �ʑA�<���A�ƌ2�N���%�ڟX��1�C(7�I�7�.^C`�1a�1ۦM}?�^�H��}mⰾ��Ô�P�d��z�Ā�
�����L@L���sx©\�� .�|�O8�g�p|?���>�)�Pr�ʗ�铱yy
��%O�w���f�����|�9�M�бZ��S��7�S;l��.����^*3�5j*���U�JJ_���46��;��oX�SА�7}���?���&������:+�^3ރu���$���+�c<���8$��n��,�J&i��\������c�S֬^�V�=&�f�u��o����/�Z�R))������U`O,'Dc�}4;��VpPRL��ߞ��f)o~�C�0�0
������0�T؋�,:8���Á0���;�OިG��c�Ol�[.�|bX��~�zzra�rEQ.�}�W.07�Gl��ְ�?�{��� ��xO>@ȏ�c�Jf��b ���+ء�g]yW!F�%9}�=%��c��+K���Ϝ�����9�.p�qh&[�z�ސ�5�VZ�jc�}�Ke� 4���Oq1����\!���I�FhP���I�� ��h�%������jG\~�_�z�ŗ\��=��&N�S�_y�v�c/��P}��W�a`ja{3?1[��#�<*(y��ؿ�����%�I���<�`�@'g͚�@>L5�#��F�^��1�`A.���ųY�C��|�� �7�����pјo�s�k�.����������O�v�q��o�;�����Y/��X���
:�%Y�d+ ���"On�<���qز�\C���?�?Z�h� ��� R ���9w�DҮd�)��:_O?���͘��}��`=�||���=O��#� �`�3��HU�6w��O���X���8����钂C,`��Y�</�{�_�Ťe����=�ዑ�a�3#�k���LPқ�2��.3.o}u{��i<D��Bs���t�<�m֍�:���c�f�2 /����\��szn�
ݵx�*}���.]v�;����^����O�G�L��T]����w��P%��l4 /���,r�&�0?�H�͐7օ c�kƌ
��#���w�uW p��6b0W��3�fԮg3`�o"���cH �9������Y�p�c�S:�_���uDH�md�� 4���o9JG��Z�t�{� �X)�rc%�o[d�8�@���.=�oߏ�8��E9��(��Ua�U�e|�M7�ϓ�yIa��03a�>�eg�������J=����y����?+���V�\��k�aa�Nv1��9M�����#�ir�O�Y�Ȍ	c#135h�l֬8��oJq8�L��w���7��>���9�q7w�~t� l&N�!��Y�S�b`��@a����j�fo����6��9�#m�� �������)�I�ce��ιD/�[:C1᜖/[�;�r���^��Vt��gjC!��������SWW���˴�A�+�e��9� ��I55)���E��ǃ�K�/�����
� w�_���<x`�?���y�I���FF�����t��4�����>#���;���f�s�7^0s�̱ˎ &�Æ�wf6�=��OkK��e:٫v�NG�F��k���\��6���n����R�!�3tP�+�TK;��#�p���*��=��u�-����}H�'O8Y L&N�m�?��{�u�&��Q��)T�7i�ҪN�s��;�Tm��N[&;b��M�[�|%����o:Oxs'���u#�Y��8�O#���I�m�q�5f�CńcY86�g�0��O��z9�K��m����7֛8�����/�F�����\됆C^���q���G�����M`םv1 0p���} ��h�.��p�ւ��+V�+�~I�r���}��Ӗ�<VM�eut�����Z��_S��	S�U���,�ǩQφR�6.��4U��m��c�]j|�f��/�8x�dE�u {�Ћ�>{�t4v����"xl~�z�9k�!���b�.19��d�{��7�o�AxʚUw��&�-���}5��4k}�:��N:�-o���3��E�⣋�披EpD�)=Gp�!:��3�;wnȂ`Cq��|�ɧ�ӟ�tp�H�p+�I�r��0�es� ҡwh�6���ӻ\'e��W�ӏw��9�T&�٬Z&	\͙�A�{)�gQ�:���ູ�	�q{af�N���� h ��w�@g]2�3�t@����e6i����~�C#�g86S�-��Ôx�/~����Mq�3o��
d��q,�m�;��o0C~�g��]j>�����=\u���𙋔6%,�nݚQ�0�E�s�����+�>G�N;^��z����Fmmؘ��5%e���/��T��X�J99�֍�a�.eI���O|�t	9��w�������B����c����c�l��Ϙ�a���Y!�l쩠���F����r����d�)f���RO��CY6�N����k�����;�J��7T �Ӗ����i�v־�N�0��(尢�` �Ap�k����i#f�qY�$��u�[Hb�(6��=�"V���cΓ[�0O�֮c�KY�|M���6�j��N}��VwWC���ҬZ��Sg�����G<����H`�%��t��"�}��w!%��x;퉶��f��JG�'�}L,�cc���ص
,�F`K�{O�7^ȏ�]�!@ ���3���6
���33�o�_g
��.�E�c��$F{ i�0�z�F�s�{�k���X����>o
��b[��1̗ԁ�A�ٌ��|^���e�F(�_�k��x���d�IH!,�LP��I���V4i�����!��d���,+bۤ��xi3&�Z04ȋ�g���%F�c��� �C=4Md�z!�qhgz!_�1��p�����0�_,X�1a�&�_�#̄a� av�UJUm�������w���	a�Pv��k7�OO���"[�j�&�$��L���7�'��d��n��"A�ܩ_�Ǐ���uji&e�'1�f=����8�jU���ե9'�����;}�e�-�?���:-9"_� �d��;2f�G�v㝞�1���=:D�p�ͨ�<Zy�G&6��
&,��o�Hy,#/�!?��b��1Nڊ�a��nב���gB�v�����6�@�#��i�`����y�Á�#O=�yµZ��Ld} '�Kjd8ȳI��6���4~�P��y����F]��a2$�!�D(�Fǲ t٬;G�;r�%B�����i�����'�`E~ ��s������l.�8��
�x��ⅹL&�ʂ��p���f�	s�'�lM`�J�w��p�*I�C���� jf΄$��F�q��V��8�Y�cA{Ų�U�B%�Z�[��U.7)�oQ��S��B�Rk�z�f̜�l8i#Y���{F;����GNL�H��zB���8��8�h�06ncNXw�'���X�F�n�J�C��M`�Lf�D�5XY�&=�3ș�%�IL�Ek@� I��A�n{�6�a�� Mϓ��� �/`��C�m�	���%?�qzz��}�=�\ߡI��U+�(ñaY�T!\פ\�5��q:;�7̽z���0���f�p=��|@�= (�A&��K"��9|�3����f!#dF!3���⸱�o&< ��]s�5�9��~�m��#�c��<�1��Yi�K�"����PP*�:l�	%wƅ]���}V����|��SO����5���W_O.�P�\��+e劍~�s�Nꡪ�T8�O���0<n(#��$wZ��*��s=Gۯx>�	0������*�0ڶ�~����	�X����X��۸=��i�=�x���quH���L(�{7 Y8��3&�K0�a�a���c�����f@x�[Lyi~fٳ�����b�Z��U��J���y�T�*[��n;k���z�31�$�!��/��!/���CQ&�$���ymo	9y+�=a�4��������2r�VlD���=�=�rc��o��׭Y�^�=b8&#LO>[y�+�1���H�z>� ̖�.���0���v���K�A>V�F��J�[?�����g4���<M�d��_�bq��J5�
 <�Wف�ԯv���)!gLw�,�r�b��X����)�Ϫ?���c`L��~k�wS@�w,ް��q���F/�ŋ>gB��8��	n�Π����]_<�u�>�B&�P�<�������;�._�ܨ%�̼v�)6Ȏb�˟5�{zU����o���&�+����/���=�~���q� ��,�}��I=��2����EM�1����X.C��-�{�<��X/N�����j��L���P�1�k�\.��k���1e��׼����7��0[Io�$4 ���%3;���@���Yn<��3:O,Ѐ�������ꓢ�#�F���zC%��S�}D-���>E�>ݡ/����    IDATJ��y�W����5�a�����CHt�3����"p�PL��6�CyE[
�ai�	ב�t�K�c�����0D��`��&k�svv�x	��p��U�gx��Yxy>���x�;�`�}�'��X���W�?��7� ��8cǼ ������M��,��dɬs(���ҥ���۔���ڒ��Kޥc��3�l��H��/��Tn����q��T3�e[�� �/�^aQ�� ��`�l��cꐏA��3 �X;]��}޸C�A�`���M8r�ܿ]s�5�" �V�=�U��1�d�cR�Ó�V4IKv���`�.XZ�ce@x�u�Q@��;Pp��k; �"Ύx��������zVi��NRKKU}�u�x�����is/ToO�JՂ
MI���S�j���+��&�{^�1a�U��� @�:f]6�1��R����s�����>�$�[9V`<��3@ ��������	O ��kv�N��]XK������1R�.���j�T���g"//�J 0l��Y�">̵,���!���{��_B�rZ��y}�/*��Qss����<�:�8�8�F�e'��?��ϭS_9���I��,+�mW���z%�}�=x�v���]�*\����c��A<�D^�C�\���z/�ǀ�^�0y���^�ך<nc���l���]t�n۽����K ��J��Ϻ
���՗\[O�TS�x0cv�'pz���y��E̼�!\����f��ٹ'hF�u��O�-�f��:􈽴��U���:����vMF�ZS�X�f�</l��e9$���M��1 �S��
��-��0>��/v���r�7�o1�<����I����c�����h����z���AO`������ ���y&>�矋T1o � �k?��={y���e ��s aV���qX�g��1>���%�>�&�՞�e�� �r�*�~ۗT��W{[Y��;4��7�ؔQ��^������|Z�F��^��]�ϵ�\��X����~6����#[ד�m��蓳Bb05��`�޲u���!�� Ӎc��t��+
�ۮZyW{�/0a�3I�0��3�cf��'��	Sw�k<��'���v���oTQ3x�%�8C}]r�{��������U�/=' �SOn�;Ϟ���R.	�d�Y�}���"Ȏ0�e<6d�ԯK+��(��`4���c,��cθ�~@hF2�c7�^�3�T[2q��1��粓
0!�ҋ��V��d�� J��H����� ����Ʊy�c����r��llr�E���DV�1X��X�c�5^$%"a��8&�iC�ӳO-ӽwߩr�[���v�	�J�O���[�U������aG�H�}��vI!�I_8���k,��	Wz�ƞw�k���C#q8��3����r1�dan0�0L�l�\O�v����t�A��wbS f&�8��<ǩ&���	��H.���C�/�ȫћ��_��~��������w߽�rEI'�:G}�mR�5T|���'���f��ˊ��qrR�; ;����d'�V�t��bH�hDf�V��P 3b�,�|�&쉵5r�{	y���[�E�����D.�8}�3>�6���͡��A/$�� /y� �]rX4��&%�6�� p�(`� !lݛ�_5�L{�U2�rZ�r����ڰq�&���kߧSN>>��-�����2�膅�=����4��3�'dP4B�D� �Y�Fr,�'��=`���A�u ��M��rp�����.}磌�:oLO�skW��^�ga.�?c&�UR;!m=���غѱ8�.fR�	��|}�J������
<��0�E�;�Zx�U��#�W넒�|�Bx��z��:������)�[��S�N'�r�^7� ֆ2��D�)��L�?�{~6l�9�W�c���C�n�l ��Ӌ�2 |f#�1�.���a��O��X����������C����0;�`�;��da��o&?!<@�����=���;@����p�����l$!E�8mlH}dǨrz���oܫ��U�<��˯�K�4�Xm���/�F��2���?�j��?a�J�^U�%������4��Ĺ�c�A�n�����>�(�XZw�=��c]6��׫����1a�-OzaL�s/G�Y���Asw ��y�o
��~9��-��CV�pލ��x#?�e`]/�s]�n��Z=��O�������ߠ=��K��a��>����ʩ��4��P;��SN���,Ւ����WyQw��^�0X��D+}<�caP�X]���+q4C�#f��9O,_?�e���;E&L���a��S����v<�� U��,�x�Ӽ!�qd�7��4%�IZ&�)��8�J�:�@jZ�g+&!6O�>�\�l����E��|^�ƕt��h֬7���G7��	O���>���w����\PWOg�?C�B!�$���nCb�6q�o8=2�ݔ��a3/��ld��%��t��\�y�r��.\���1-e9����x��r�aÁ0�����]��c�A72�'��C����5�\�x��B���3�v�i/�	�n!1�Z���?z�j�U:�o�g��V�g�u�POOa �{>����C����B��"3�E!t<����d�Z������G��ً�+�|�p����Y�B�	�`FmX,����E���/�]�>��t�� ��<p��ɒ��]�B�qo�u���v�����'ǁ�qg5��|aT��w���s�m��oPss����b�|��d������?ޭ��Ї/�V�f�l�(4)�M�- L�i�6<V��i�I@�8{����vl�z�U̃o/\��}cz�F8����{u:V�'LL�ě5L�T3b3��:0T�'�n�y��<���B�e�|O��pD:&��S��>��oi��:�35uj��{���ɲ�<=b�N"��#V�'�3�z&��11f��&�P�nk@m$�{Dą�o'��<��f��'N.[���]b�.a��a����~r�d�m3�r��a@��7�:�d���=�F�v��]�)� 2� �yƄ#	��|��9D��C
��.yN��M�z��Œ���/u�)Ǉm���=��J=��J��4�����96rp"M���|���a�� �##�����66����8��a;�wa*/�zm���#�s�ܷ������9�~�u���!#�0����
��������B���=1���-O��@`B���cP6X�r�7����8;�q�
ɰR�Q�nפ�vjҋ�*��W[�6z���:�����ʐm��:��5t��yz��
��$=-)$���y,�x��A�1 !�ȴ���X��.��G����?ވ3�V۸C�gs�֦&?�u.�=�V�3�+�b�Q�7Ġ�^F�x����D_��ec
�dl���8LF�_�%|P.�n�;�q�pQ߂����K��2��@�*��زH�khժ����I�r�&L(꣗��S�E�:E�
ji��Ξ��[�J�FA�-����W1?Q�|�*��"���\wi|���3��u�{\�1��I���PQ���qaH�C$�W= �ߢ��A�����M��|��g��eԎ8� ��q5�#��~Ǡp�Ր^cpuz���t����W�bBL�=�0�p�����3�(ꌠ��Y�����7[4O9�A���a�TQ&ӭ^xF�dU�_�b�-Z�lI7��yuvV���T�t�����9� e-I�ګ���|c6ʢ'qa&w� ��cm� 	�2i0Ƹ�^�J�Gb�ǵ%�&�W���'�}<�@X�� �	@;Ǖ~`��k���o�8�.�@�g��u���ʞ!l���dC�>�o��!D|V��Yo�c#~�K!�Ax��%�p������>�zӛ�T�ҝę�ֲͪjm��b�8���a3T���ib�I�=�$�h��6'�5�c0�G6)��qp(Ƭ�G�a����wv�;��s�yޥ�N~q�ɍ��=�]a�!�J�,RԪ��fL����>v�hs\T3$ǁ�������Xx
�s=�q�|��'�|������S��T�{����˘�(G����xw��(mz2�uU+�����]}}T���">�RC�R�::9i�|�lO؜2w��|�5a��$�$[�_�?��qYD����4��e�͌f4rQ���opӃKY�
e#`#k�7�`$wכ,�61��G�"�!�`١�a!l��6sX;��l�� SH��������~y����Z:r���;�YI^�p���"}�Q6TQ[�b�����HU�!7�6�O�m_ԥF&�RoQ�ﰫf��&L����B�����dיK�z��c0b����7��x�	�S�X�d��xa�s�%�����H�Er��k��g�End��0�T@�Z`��{3coj����L&�\8�Lxƅ�m�v����(`^�6�s�zM�BU3^��������>!� �ԧ)�H�Bh6�Bz�:��@3�u��t>��yw�q��������PV~��o�&�0�c�9F���g^v�	�cZi�|��!$�У�>�Ro�����^M?I=]R�i�*UJ5�l_X��{�ٚ6m����X쓣�^�?6`���DQ`�;p���w��h�³�*�(�C"f��-�4@��|4��^ރ�xLlBo,|yK7zM��v`��d�9�� ��3���f `��9 �x<��x����`D�`ڃ�nX<�ט�,}��{:2�#�>�;ݭJ_�*�t��U����q�p|Q.7A�}d*�IS&�yCK�=�s�0�I�tE4�O��	�����a̚����� s��� �k��
+�'�`�]�ݞ��u��`$�4���K8 f,h+����˵�^{ј���,j/��p��b�®{����6�Ӳe+B���h�M�K�@�J"4�]g��5 ľ��m�Q�N8!��}�����gs��fፓ5p�-#�;��#f��3U�to���K����~�Ҫի7j¤mU�g9S$Z@x��P|>O�N�}u�178%(�A���j}�������|� �DcB�v4�Ǡ�c��Z��L�/nͻ�r��8%履�#�it]d���iz�d���M�H��C�`��9o� 0I�7��p����w�6��� �P>r�^.�X'�����%����kɲ't��U�mRS��\�W�ҋ��-�*�m����@esM��	ƫ^�"bF�}�P:Y�\�+��8:��@��tµ��r�[�s�}�7�ac���H,3��ZF�6�`��]�1K�����1�e�Y@��c��_�hۜ"��<N�jV��m:a�����{��?@ؕ��xfE^0�$!4�±���㸕'2�b���s���(�u�]����x�_+������ٸofo1��چ�*�6�_�s�:7vJ�����sEe�mz��U��[U�$i4� <}/��Ձ*jM��R&l�4�dl��3�2X�<�1ak@o�{̬�Έ�7���x�I@0���ۣn�;�>�X0�	�9�H��l	t�z�|a����:˖���?�i Y� �ș�p-2�~�=�;w�0�F�VM�
��f��UH/��?����5�vJ�JI;�8A-�R&�d0��8q;�|���m�}T�'������{�9R[ɰ���y1�~;���81���w������'�3�� ֐5� ����*{��g�l�����³����p�C��[�^��r�o.X��c�SV�^4%S �i��9c�~�5�Z�f��z�i��&�B�*!�3�!�V\��N��� �^���{Ă�"�&9K�$.��<�����o���ͼl�`�����o�)_�R6ӣ	��U-w�����{d�.��@�	��4��>��|~@yY�|��YO�f �ǘ$� ?('���΍�lDc��g��@G�0,���Ys��Ѿ{S���KX��3�&��	�sl֠�.X3���C��i���y �s\�g��\W��0b��;�U��)�#1��K��60�'�zT_���j��j*J�;O�f�\�B�v���ꮄ�����h��ev�����)��2����A��L��+d�gȒ�:�$ ���y>��@,���:gW�5��N��^̴�y>�s �{�'`��Q�V�����r�!��D�6��pso�A�����+�SN����_��~ul������r��s�(��M����(X���ٚ̝o�2���!��8���dG���e�	i_Ҷn)�N�nۢ���ɒ;ث���z��:y�{��פ��j �,���|.�W���dDff+�9ed�����-��a�5�y���5�d,y?���y�=*��h�vS�g�qYЁ�B�K��d3��j��/בֆ�9����@�(I��x�f�qxs0�����s�s�E>/p&��49�Zn��g2";��/Q�>M�ׂ�.Ҽ�OT��Rؚ[����auu���P�S����d�l O�s�v�X!/�
#�#p��=a�#�u�r�l����N
�x3�מxD��.��&����7^�䏐���Z�V���},�xLA��)/>������B1�r��ݷ�U�z�;�b�Z=���b�1~i1��Sh��`k'?v]qP*,44�ů��\���Ș �����Ზ��<I�܊��X� n�У�~����L�)sߢq���j�ji���U�o��j ab�a��K��pD±��@�UL>����B��N���l<]d�c�:���3y�R��}���� ���@!䙢��a������:�݇��aa��88�y.a<FdͶh{0~;B��q ����Hy�=���l���m>�b����/�V����u}貳5{����e���o~L<�f�8R�l���
;�Z!�̚
�E�O��zǜ�l,[���!�����!��v�w�y��w�yg��E1�1�d�<`������_��R�����{'��"]]�֢j�|���^���1�k�/������NJ=h�:�y���%O�t�#�0�!�Kh�]4&�Y�Wym� �\-r��c�y����F� /l��o��E��{b�P�L8��V�z�_=�kt�՗��g�N>�X]����5�G���y���E5��x0�/��9]Ӧ�|XGxɅ{��0�J�Γ�c��;��Ŵ�ٶdru�W��Qy�x�:���nh/`mjG�h�e�r�����β��i`�,�՘�S�(�ü��0�a8.i�-�0a�8���c���N:d�35�����d���Z|םa����U}�w�3���?y@��?j���.�kM�v��բ��%�^V6Ǯ��td������aLa���1�<�G�Kb�,ԓ����O�!ț�8)�5�9��)������Ż��l/�﹖�ID t��3ٺ_��j�|��kn������o���ֈ�5&�Z�hJ�q ��t�̃C8��?�ZK�?'��BH�0�
���;n��P����.��� ��[ɉ��x�A�l�@ ���g�pPZ��������p/��@���(p`x����_.�u�]���zXS��붯��^��nz��:�B�F�\K�u��9�����d�k>ʓ5�I`��} ���zP���Xm̈�DF{-�i��88�?�b<��{<�}�A�߱[�^�L�O�����[��v/��3& O�u�sp~�Cc|�gH�&�5`���x����yq=�0��L�|���-c/�� ��X�hb����V��oUϋ�0���^�N�|ʛ��]�5�������4i����G�����U.OvUF�ZU�BN�P'Y셩k�I����J������Z�#;X��?��p�����xA��~ثpx�ޅ�:��K���݌	�;2��}q���E��W]=L����~h�I�W�9��H�VUԎ8�0�t�,���/�n�ZUJ֓�5X,2|2�����ut
A9�������v�m�s^q�3 �-oyK h,��,>���0g���_�u��9vcE�qa�sl���S��c}�n��:=��o5~RC7�C:��Ѿ�q5    IDAT�uݚ5���4����Z�"'���	�MQshd(F2�Lw����l(��y�E]|��~;��+06��\��㉀m�B��G�V�5}��I�3�aY��x?� 8��6Z�M�v�g���.f�<P%��� ���qȇ��0ۀ�� �2�ŋ�[�+᧟Z��~�N�z7h�Ć.��,�tқ�am�.��=���~�}��_��4S��b}	0��/���<�f]���g��n�A.0�P��s�f, Ɛ1Ǔ�]���3�y��X��;�;9���	��������6!W�AX�b��֔����]~��z��m[�#֯�����P�Y�����ЬYoӯ��־�F}=����D��d�B�,OPB,�58l����ɂa��
�����{  ��Ib��(��t=a�3a/,�)�ro�nXx�~�˟��Cv�?|�Z�v�]�?,�9�H��Y5���
�e�� z@���F�1�RR�g��P�?i��f��<�q���s�ꭝd�N߁�X >c��ǘ�۬�qf���f&���K_gC��5{"�`e=�6
�k�x>���c��aWN��"`0��.�,�9�3�7�^�Mf��K�¥��\sD���"+��a�n��~���+��[յ�M����׼S�g�Ύ�n�����>���t�?�LW��)�Y�(�YQ!�{��Oh�e�¬R����w�;�l�r�3�����_���s`��#L�x6^��+��m����Q�QJ��"�E8��R�T-�͎=����ի�l+��R�QML�p��5K��G~7��!�����e�QB6g�BƲ $���_���+�8��ěY���e�vBA�4��+�NU�~��>�7k�LC}]���+�ѹLg��D��]�B�ӧ�\�s���[WW#ۢz-�l�%���
l	0��9�h���Ō��,�-�}a���e�¦fh�@����� l���^�ݢٟ�x8o�+��8�c�h����6Hq�G���{ ���g�5.$c��
=��X@c����3/�CΗ'���x�KtP�}{�<q���sk@���+���;Gtj|{EW]��r��[�������S;3�����}�6>I'$5�yT#S*I5$!T�_W:s�~�h3��
���"}�c҇�c�`��@5A�x+`?f�� /d�����H[�$Ƙ��?���z��"u�\u��fG����z�0����^����[&6���ab���7����<�(n�­ fC$.�LV%�w�:�zK"ʉb��0���IlwvĐ1�lM��F=��/��n�5c�.j���J���/��Yg\���&�5esy͞}�f�<0� �誨�Y�A��O6O���dw�w������k6N�b@J�S��H����i��h(�m�=�Ѽ�F����1� ��?��\�F�UG:/0D� �\m���p���w�AR���zb� p8A��G�M���#��Kw��ԳO讯.��\����L�r���e��k�~=��M�fg5�L
�*��Z��ve�lEO@�m��$-;"��q���n��"�	P�Ff�;l� 6�,R�LҐ��W��8��s#§n߃AMy8����1jGd��o\;�y�1qՊœ���j�Զ�zӛ�ӌ�����Jk_X�r9�c9E�Av�項���a��A�X*�j���b���ISC���$@���Q:3l�-�}��/+xb����j���V�.�L����׺��7��?��9���֯���mV��JnA�O>}�	'y�c�3u&���m�c �Cf�q��,4^�Ќ�6�k�׋v�o`6 ���e8��6�n_ړ�e:�$n}R?$�?cc7b��È!+Μ ~K|���`x '!�+@���6{�{��\�Y�?��p�b�̛0 �}�7�K!=��?[��.}*d'�<R̕t�U��ig�Z���T&�$�V�Xޡ	wUOO]�zN
e��jToY�<��x�7�����S"�����~7l%����L�!�a� T���K�"o��%�>1n�'�
,�X@�@��6n����������������ï������J=���1�L��M�Wo|�B��}B��	%g`mM��v\ǹx(�! ����ʧ+b�Z�LB
�\rIP0@څQ�Id��0�aet\��*�'z:~����R�Ӓ%���)�L��j�S���YU�7�����%G�$ LLx?e2ĞQ�х#b�f�]f�˓� ��.��l3�� �H��u�&�A������4 z�Gz�pߧ�f�N�73��P᝭iG����{b�3��x���a~3����N����u;���E&�8�Cx�� ��P�Dr��)����D���۾"��j�Kg�~��p�~�zT�R��MM�SU-OЄ	����������JT-l
���-s٘apDGX�!�@H��0^��g�&j�xӘ� ;��;����P�u#֙t+ި搩A���	<�ZO�����|.��k\;� �M��řkon)fX�ʔ� �qo=F�gLӒg��s�%q&�h,�`�B�3������2�ʈp�^\CHdF�
z��w�+��Au5,��7�blN%��`N��$���l�G~��֬^���^57eB"�fM���mR8����O �IQ��ד�)UN�3c
pܯ��-����l�l�=q�y�-\1�؜��k�kE����������h͜<C��t��c������
g1�m���/\�3`d>8������8v�wZVl�^���m?�c�2���z5iG���u\U�q���	z�Q'��}�s�������|�/�-�jo���W�#�X|���h����îC�+��G?�YT��a0���q��
u���i!��~�7 �aT���F.��Ƃ�_&<y��w6uo<&�Ԅ�i��l��O�*��]�b�։N؂��C[r�e,
�c(B'��vĖ�g��F ��=B5�5k��G���␄]A��1c�|*K��/�鬫Q�(�k���Y�WooWOR�2�d
�,��Ve0����&��هc��,��@y��o�'^��A(aČΟ{1y�/�,;������K �1�JV L�P����F `�O?�ϙ;��Pf�\k���/f[3�	��e�t�w�^Ω�H!��IA��6�z-��	���λ*_�T�q!Lx/��7��$Ԓ,&����|N��?��C���� C�ϟ���7�8���>��]���ο�R&cY����Nj ��󦒚��s�V�5�-_4���V,n���/d3l[v=�Z������POx��v�c>N���q,��1+�)����)1+����b���w�3�����Rc*y��6�%`pI�q�%��%1SE0��>�J?uA����
;x
M�/T	���Y��e4w�;4m�tr�Qݛ�~c�d�n]ş��nc���$�g�y"�8�~����������@<;�=5��F �����t��t{�S��g2\�m�G���� �t�R�v�"���.���p�Q���zN�B�z��!U���M���ڦJ��l�d�0�6'ٛ��x�,!�]���*��n;��a�=~0��y�w�DMa����xC�C����O�&^a�\�r �X�`�+�m� �dGP�'��ic�z�
Y�f���Î�34����+j! ӫ�\� (���z��ư30l� ��F�\�s���t��H�Â��f��_�������~WϯZ�lnɅ�Z�z�	�k��+��g4m�~*d�����3�<)=����%���qB[e�E�i�,��ʭ���{��i�|����x-ē��[k{w|�%�7Vc���U�v��QS�ګ�v,h�m�T������є)��cުw�C==���A�b����?��N��$d���u��s�v
X�6`^�3`6[�lp2��,�9�����kh�: l��^t�=�1u�w6uw�*jo�7z��ʚ2e�`]���mÎ	z�#P�2�Kl�;Wb��5a�7qa �;e��c��x1�v��n���r�AZY9c�^ߠb�������.��j�z������h��5��B���@8�����[2	�p�7�xW����t�3��dY���n��|�pO�������:	�^�	Cz!6}M����Gb�[�җ�
����������ޖ�{�{�f�~��>1C8Y�V�m4�IjK�I�ĳ�����m�x��/,@�M+�i�r��y�� ˜!��6b���g�p��3�#�Q<_�y6�\6��k�9މ������"�1?Y� ���yD���~Rq�"��gB5��`9X��2�@30�
O�1+-�5`L�^��B��Ya�X�W�z`�@�X(א��A�q��j��B�G--%m�C�
�%��_Tk�=�h�N�w��:��6� a�{���-�� ;�)F|n��q`/��13Jjz1�qrRr,� ?�	���o��1��� �e���L�8���[ߺ��4�|�Y}�+�%�|����/t�;NPw����W�>A�W�k�z��q�_X8�r��y�>��Ǝ9�c��U �f���F�����-��]�q�٤Ћn�1�@��;�I&;�:xŏ�׸�QL|��u�]7�g̑�6>"��5)[&h� �!}lZ(��8o��6Q�v�*fet� �n�]�C�>f̎�2�����ư�gN�I�A�����ߣ�v��c�?D�'��W��%%�q����*��� �p�ys�־�NW~+@��:�	����)1hDS~����7�12�j�1&�+��gZ���u�1�t����X&���Z��}�/�V*�������9��R�K�B�~��r���g5c�#��v{�^o��J�.��pZ)j<&�s&f�7h��Ldg�6�ۺm�p?P��8��Ƅ���B62��z0���]����F�]w�y? �㫥#�1;&Wj�c�=��8�<V�8��t&[*���3��}�N*O�6���1U�����S�A�v 뵒�}��Q_�����t�E�PlҳOm�ɧ�'��Y��Xb�[�^���:{[��e���Id���v_L3�X�̴=F���Gh����J��h�����C��بZO�γ��T�q���;��Wb���K�<���z���;5eJN�~�l�r�q*�K�����>v��Փ�G?z�f�<T�2R� 5�pO� �d�v����������Ƅ�ޞ�c5�r�5evmF�8�1�އÞ��S�����n�a���O�x~q{�/�0g���#��bU=9,�Vāp�q+F�:;ǒ� �w�xq΂��f oK���ټ�L�85 ��1~���V�ʽ������k��L�?|�cz�k_��˻4��w��/�Z8�4�rν�[.~iFb�ܰ1����w�(��!��x�c`��bO����Г�x��	$6��+1����Oa�e����x^��X�����4����X�z�]��٧���ޣ���v�5i��iμ��S�u�~B?���i��]4���{����2A��^g�_�<,5�qK�����):�T33]�nM@Lr�W/��egP������+^5��>�ûW�/��2��|�n���X�%sj���x���'�yaq[����ld�����+�����]c�Ke`J�Y��mS��O+v4������|f�EV�~q�>��k�裿R�(}��u��k��>���3T�4��9r��	N�7ڼ�5�@��̀��`�El�����ld����D����X��(9��]CV��Ɔ�-v�F!fk���EX?ӆ#V�4��;^��3#{Kq�ʆ����3���I��x��A�Y�����8�kƽ���i_3;��`{,c���X���G��sZ�d���vU�]�0��_v�N�}�:6v���\���
m��>��ŗ�W��-iܸ� �l�pQw�0;x��զ�U���Fh�~m���Id�\{%�����#BRvt�m�.�4�7wЇ��wY�Vΐ ��|����{��K^�G�_{﻽��Wk���ԓ���i���R? \�	�dan3JY����q�B�Vi��̛,T���꘻��1���d�=��1�1�z�!FݴR�3��Y|<��p���%6i#3��6ǋ7i���5����-�L�c�g�n����ux��������Põ'f���G[z����%��J����t���ּ�NPWW�>��O�ޯ=��^���ϿR{�}@8���4N� $AMn�W��u���A�����i����:�����%�S��M���'��^:�o8�jaœ4�vK���{�b���S̄c dW�po�.��|��kt�st��ǫPl����Yg_���A�>m&<��s� 3A�v�?n3���bOz����eo�@i���ǆi�g 6%��@�`�4;����wm,�GiZ/�&����u�q��:.���ٰ�š����H��c���4�r׻<"m�Y����f�Eǲ�Y��ѭ�W#ݗ�OCK�-��E�T�/������Ь�oP>W��zH���۵�#��|讀1�p�Q�?���4��$���s��z�`�n$|����0�Ɵ�=��0؀f���&��f��N�'�[��:9�Տ;�g�Q�qU�+aO������~��ϴ��4󀝕-t�l�������Q�:Y��,���ԱH���1� �l>�<.�9�k�� b��y���n=��o�(bvf٥�ᦔ5f�1�ĉ��i��������b&2T;�No�u��Y�~Y�}y="�$�%RiO��c٧��,6�d�I�e������D��!3����1��Z�sҞdl��bj[<��� �|ų����]Մ�y]qջ��YGhܸ�J��V���������M���z{)yYT6_V�ZQ��2�$�K_�� � l����H�X�{�P���5��_�翢 ���r��ń�pD�CVʴ0��ck���1����Daa��V�� \��Զ۶i�]�iC�RU���6^O=�^�x�ձ����/�0�-��>�p��@L|( 5Xx"yU��{贗X>�Ryp���'!���s��k�a?s�v��4��[����e���������:o����>�}�����C�q�؀�k�f�#M����^����Z>������>���Ǜ�x�J���,3��3����� �ٚ��x6�`�Y����>��$E-_(�T�	�w���=ڰ��9Wrr�1���#Y)S+)��6�H�9ֵ�H�H���M��Ga6kLY�zq[����@��t�l�(�$i �d�=#	j���<610��M�tJ�����U���d��Śr�>���[�yd�>��E�x�z��ԏhd5w��6mor��c��L�>�x�P�|S���p���"fαu
�Gb��.i���ń3��3hx �gg`����(1�1�4����)�!p��2`{\b6��}p8Ǚ9��a�5�vJ�A�v �Ά�����:�a挌Y�w���<֩��7��/�W��'�I΅���4i�8͝������Z�̙J�) oK�d��m�f�LQS���J���`��{ｃ�ͦ͞�B�)�wsI�����ޡ�<_w�u�t�Acw�\r�|z��FCeGp�=B�W���c�.���IY<!͔�(����Rw������a�������h�굡�i>WRSsQM-mZ�zcP�z��l]n�5wΙ�6}/re)�	dN_E-f/���7{��pb���}��J3]?�{CM�l}�(i��B�H(Ļ�x�����c���H�����H�7���oo5EnT�Q�:v7�vV���En0v ���N)C�.��i��R@�<Q��=���cEǸ�]����x`���Q����Cޜ�g\�ߴ��
��g�����/*��e�i����	7�b��PO���,5*�8��bSC��^�s�j�U-��:�����k�T���G��H�.��L(?��J���P�O�k��M�{S >�}t�s��B���	Xx�x���E����\6�"@t    IDAT �< .9�03-����SY�z��.yF]��SsSC}}��+W4q�d��Sn���
R�0�����~e�y L��2��� �!�%Č(�$b�|c@
h,���D�aƘ]��9f�~����� "��ras���K��ٟ�/n k�a!ŏ����8�m��|츞�r?p@���� %bx�Ϻݱ��?:D�U =�x�ϊNS��
8s���T���=��C������9I�q�Ɗ���U��<����̌�p��b8oh,w�g% �U�G�r_+��^ݠ��L�I[��TTSk���k5QV��ZhVo/ۍ��q�^�t8�ۃ1>>�}86����M��?��I�qɺ����@8��|���ߘ2a��<��([��B�0���I9A��A�cX
�,�5NQ<��}�׊D�< L^��{�A0����MM	&ŭb���[�1P��(�ٷީ���ڸ�O�Ţ
�R-�\�k\���ԝN��>���S�<R=a�>���A���4x[�.��Z�(iV�sm �ﲑ�Ԅ�a�Y�}1���s�x> F�*��� |�nP��ǹ_���:����� � ���\Y�y�S-p�sJR ���͐�5�w��FJa*ڈs�1l�g��ϸ����������h���Av(�� ������ (T�s"0流��G���m=�n��A3=��3!E����^eգr��9�/kVo_C��O�{�|s�j���M}�l�h�:�3#����/�)�<m���m`��L�^`���p�=2�Tb�|"	��=�^'��z��#�q���4PO���^{�؂���~h�Wߙ�XHKk�jՆ��ݣF��LN�����S�冝�1�E-BA��ꔫ�4%��A�if�Ii��I���B��̘1#��b ����G�v��@>_U�����[]{B�x�����>Y�>�<��7�I9�F1	GL�'�!&A�ˑ@0�2������l �FG�A)��Åtb�3[��5�$	�1�iv�{�:�|���L$�0��z�{ܟx�ĕ������R|�S�gr�����< 퀅`L0t�{�Q��Xo����C��<z	�@��u�6�S ��)�އz(lЁ���^@Ma�C�e��w�>���;E���.^�zU�����Q��K;m?NMM5��!&\�6i��u��ў�LW�RV�*e�.Ԝ
�$�P�` t/��2��#��b�9c@�c\���!��˸!_��(Rp=0�3���f�:��y�K�w#�����W_}��u��#�Lza٢���C�[���+�3�X����*j{�fO|�!m���Aa�f`e�H�d��Ը�>��;�4����5��E8������B���/|!���$�bya�@d��Z@�)_R��1�1ǙX�b5��<��]r�U��ͪJ��=X�=�1����ܟ� \��u�Pc����,���3��k��r�,>��y�G��	3�6�����0^�������� ,�8��(������\�������N1�0
�t�	0ia�0�ab9��w0�i���|Ǆg�>����y>���  @9 ���+���Q�T^�I��6��x �@tC»!����4�q�Y���[�C��p��O=�{�v�*}M�Ь�Ν�N<R���pe.ӦR�E����o_(��VON�A/���`��?��3/��<)g��7�9��c]5/��60Y�������1cl�27T=a��������{ǫ���l@���\sͅc
�3ϻt��/�\4�^9�R-)�ɫ�WSKKs �=�z��>������lM��lN�q>�7��(��Q� 1
- JO=arsY�Eh��T����[B�O������}3��,ۮ���T�8�+���o���M����i���R�@��Cج1�lM�w?�s0��A�ﵑ`���i �;� f��p^��ű������8��V�,�@76ʐ��bHc��Hߨhq��k]q���' $��K��γ�O�-z�'N��st�I�u���Ћ@��v�Oȋv�=��a��-�����29ai > ��_�@�0l�5,��q0��C���v���^r���0
��c�6Ң�Xo���z���s�"u��P{kNW]�>�=��z±�-�m��ڲ�{Z��YW&۬j� :l��K��.�{���M7�<��|�;�O<��`h���y��o�G���u�܏9�0n�/޸��r5�r<�x������"G�����n�馋��o��["�M֎ ��ٰzQ[����R���&���N����4Y�Oy���v=��s���,9�f}�a���Ą�pf��~����N�q,��p�
��<(?J}�y�k�UB�?�Ov,k�<x��y�Vؘ�e35U�6��?���ݮIo��Mݶ5���S�:�̋�ݕS�)�� ��i���*�bx1����
�X�Ǳ\�t�i��q
�9�Q^�H�2R8"�	�����@p&Ɵ~�)����7s�<��\ȡxU +z���5��	��q�y}���C(��`�.��;B��"��<���c��0�	`��:>G/��LpXυu����0fX/s���,��9j<��Ah�?!�{ˑ���� �乧�h�������Iͺ��s��YG����J����f�~q�㚶�Q�i��jd
�د����F������#dƸ^q���Qo�8�s�!��NcG� ���z��y�������8��$���{�a;�������Qq�8 ���~��7`LAxƅ�Mya�����'\)�B)���6���t��o�#�TO>�t��^f�h�]U��R� E�����s0��8��f�p.'fP�߼����x?����)[�8~�������Ї�SO�
�9�x}��sU(4�G�i�T)����0y��%������B�����p��V�����E0*�a�L���c�~�A�r�ӻ�Frg��c�n&LȀ��SB7ƞ� K�i�f�q̍�1	a,��3 {�9��yc ��|H� ����[�c��41���]E���B?�D�k�m������� x'c�w��ť��0n�H���n�ﳑz% vs��x>=��i�s�W��թ�m� �s��Je�~���u��Q�:Q��M:����y@�Y�������R�$��	��� )tQQ:� R�@B�Q�qG�QGfH�
�{g�5�;cEE�����S�~�o��9��rJN`֝�u���[���{?�����u����!G%�R��e���S��e�]�!8�b�40S�Pa���I�A��ڬ�3p}m����@�/�'�6�ߋ���q�8+�J9��>z�=�\7� <nժǫt,��nڬ�u-:����w�Y��z����ٙl�G͆��X�3o�#$�iӂ`~����b
6�Z�`��0ر�! ��1U𽽬�ۢ0p���U)���5���1=����k�F}�>�IS�虧������0�#*�L��-i��Q�'�[e�=�A���o@�
m0�s��km��@�s�n���¶����{2pa~ L�Ś�0��L �Qz}�*�E?-'�況P�3A�����Y�q�#��JPl��͎K<9ޡS.�ͽm��;~g��Y�@p/ƻ��k:r�c���B6��g�s�"��+���e ̭�������K�葇����ujn,k���u�Egk��պ��껏=���?X�}t��r�r� ?t	iJb�y�<�@_��W��6p�g١���?2¼ cb@���l����y7���#ք�X��i����X�ڛc�{�k9�N�:u���Y�|̠������?�е�X���">�g�q���6U?��h���P��0����a8��cDg�Y�`2��.x���E0<�C�0@�{X�:���zo��jG`��li���;tӍ�ʕ������go�[�v������U�U������9������Y7xt�A1��	���OWA��L�׈A86G����x�̭��`7Р�	�g�s,� 6MLV��@�Ƶ�m~q�P�ν���ڒ�	/�q&��;6�p?�1cԑ���dd3�ׄ����9���Q�C/�\�~9���v	 �N{��X��皱���s+C-�C��+��+_�??�U�^���h�7|Pg���ڸ~�n�y�~�����u��kn�aG�R�$�K-�F%�s�r����!?daYǋ-���6;X</��wh�<�gd�Yg�ٓE�9���>Y��+��3���g��= �i���	L8��<r��wlXA���u+LLW���� ��艺����Ц���7!D�d���6?X@�$ L��A�N��P�PW��>еM�	�c;jB���>X��dprj*��#�*��<h��C��RG��ϿI�-�������Kws��v�<�
��Qԝ���t��P%j{KY���0�OD&p���A�,�����bu���|��!е��&llN1��J��6�x������`WM
$9����`���C�T��Y��ǹ����E���W�C�`��_	g�K�����s�Ǝ�n�s�{���U��/�;���Ə?P��Z���jsg���Ň��(���15<���}�� �L/�>�&*k���b�.����p���P��oN��^`?��o`�&���D�Y.�[�VK�l��;��������l�w&:b�����sgiźez�O�14 t\�դ�	 �ax���N
�;2o̚=�	%���k�q���� fT�/���V��t��1gGV�a�WJ*tm֜[?�be��=�T}��3B&Вڃc� ��l����9"��3��cbS��3���O
��|��a`��8���06ؔW�X�1P6Ma�m��?@4`1��ǚi��_��@����w�cb��5�Ʀ����#��tQ��;��+�e�Wj��_W�k��[*�w���5�=*:���	����В%4�_k�}�W.�U��{�|�a��::��
���%�\4.�M�Ih�?��OA1`� D�s�	6\L���ڷA�"䎨�X3�0�e,d����R.���]w�qð��W�t��+��7Wߐs's�N;�T=���kɲ�!l��au�����@��`�ǃ@ '�pBx(؃Kj�4;c�Z=��c����q�Οv�i��.��%�os���-���ҟ�����cu�Q����|OIK_�Ѭs�VG���%�)͜y~a�\���µ c 4����w��?1Ǫ��A�ks/<Vsm�����LX���ju�{8���; �m��N�Ys/�^�G�5���s{�����ׂ�`�>>vG��ζ��8��h�zh��
ɦ�7�tipp74���Ӛ��z�wK��>G��q��ne�Ⱥ���T)�T*&Yq؄!bk^x�L!bD�xnجd�/�;�gy�[���0W��=�v�����0�
3' �{�89�lF���6�';1W��b6���Mw�����&L�ܸ�5��[�'c�舷�&�z������֮_�j�B�b	:wG��xP�^1G�[�����(���
��*��w�}a�
D���g�\/o�9"�x"�S%�/k:M���&˛5z�D���M������`�% L=a2��L��]�]���� �An�!FFqh�@��L��l��M��`�Vk�����^`��MO��$f�Cɥ�����5�m�����p?�9�K�J�ٶ]y���z�٧þp�Bݕ�s���Y�P���U�~��ܬ���^�ƾ.��\����A!�����&-��5���D��BRc��m�D�x<:[��v�����2�L ��	���1�W,���}cre�nظ��rJ��o�}��ӦM�8�P;b�K���g����<��t��g�W��^Z�2�1ǖ���A���#�!�=8Z�.���Y���r�uׅ����}�J��(�m���/�� ��@�-�m_�p�Gi��mzy���Ve2y54)0��Ͼ����_�ё؂�a�C'k���>fr��D� ������13u��P�C�p��X5�Y�ꟁq��
���MW����Ү��L*;bnٕm|-�m^�jY�Z*t��Tt�������fHDO�(��yO55�r�.)ϙ��A!���=}�����`�2����n"�K�1cF0;����{��̙�����:����;�@-��B�YͿy^r<� �p9��磏>����t���΄]E���9��դ5���4s����y=�̟Ö�v��c�p��!AN�Dh��@�`��}p���#,�3+S�Y�3��6�$��1 �U�]:SQ�5������6mH���*��qcv�K/��Z��v3��؄��>s�4�J�ⳳ�~zU��E���t�9��[˫?�i��sG 8�����֪ݖG-�0��YR�:_&�� �Kj��4�������l��*vwh���ҩN)UPW���B��1z�)gj̘�T�Шb1�J)q�Y�1�ݖ�3���μ�|@dy����GG�ܘC�B2'a�c5q �դ��O�+r>�&�{�������.��JB��j���w]���V�؄x�~:��)�(����R��x���6���z�bV���P�6G�9���{:Kܟc�<�b/?̖�!(�:�q��*�h�吨x2yңN��CJj9�wu�I�L�:�Ⱦk�a"��:w�y�<���A �)q�ݸw���1�:��H��;�m~qm�y��1���w��A#��Im;�N�u0������<�%��xQL���j,���ᯠ���W.��a�L�	���\���TW?N�BZ4I�'�|1qd��5&s��^s��z��fln�{�Ø�$1K� ���;���!a�1А�B}��_��0V1� -����&#'�6�J'�!j�̷�c�Ǐ<��u;����-���=E�6jB�	�a���o~��M��c@@x8� ?�,�4�,��:�<~#�{�w��� ���Q3D�I	�A��2��y��8�!���,:�&��B�[�<��
��rlwTج�&���kR���p5�J*���,��w��D���88� b��<f��q�c/���1�m/H�2P˯���}����<����As!��ׄ�ϵ��U�Ȅ������3=�yf�����`���x��C�U�$@K��|!�l�I�N��Ɔ&�����T	W��E�x,|mj8I֠��F�4,�^��l3Z���`8�v���a�0a��!m�9���F��m�Z8!�d��l.�J�\6��=��9���W���4�	7�7��Q�q��3��G+^Z�%/,U{{bǵJl�<�l5��WNm�{-�f5C����k�C���W_�C9��%��	� ݡ-�U���1�[l��Bq�~�����I��Sg��~C�ʩ�ҙ\���3�Sʒ*jea�I����L��sF$�jI��dj�X�g�v��;锖�\�i=���w�j��G+�KJS��U�u�m�}u�1o�GLS{GQ�JJ)�WJ��i��������R��K/�4�p�l�/�	��~!H�9��)���p�{�w(h���66�Ӭ�cC&t�����ߞ;w�u��c��qkV?4���V*�:d�)�������8I�M���Ͻ�ի��q �M ����0`�}̪��V�">���������b��
�*F!l4_��8;�͌�cε���*}:C���*�4zt�Ң�h�2���x���o�jU��� ���0�r��3�Wk��gD�!�W
�.Z�@ULu]~��q�)j�˨��H�Ѫ���^Q*3Fi�V��R%ӭ\:6�����Ct��E4�B�3gN��w�D�>�8߉~ ��sX  c�.�1_��`Ä��DJ���t��Cr�Y2f�6>B    IDAT&��];Y���R��调�����	Kt;k���!��}g���l�֭��}6^Yl�WV= ����P������v�|�PҎ)�1o޼p�PGTH{��߮�|�3!J"V�$f�-Ղ���L���l�F�ɨ��U��l&=��պ䒏�u;4�
��JF�g��)��1W�R�`����pL��k�H`WH����5�������h�u=�3�ÚuJA�,�њ�Z��G�R�Z�^�|-2�����K�Z�,;����>��`������ʃ=���������!`�kӣ͛�/����Ô�(�
^8�ӱ���W 8x��_�"�@�l`�Zeg�]»mX�P�uô�� 8i��V�iJ�I���ScƌN2�÷s���8�֋3&U{,3�_�g�(�DG �ޙ��B��te�`����C�j����L�ݖ7nX�_��:���:��7)�Mj��y�K���Zs��E�% ��1�P�	�����
d��&�W
����}�+�fRjn,覛/���:Y�9�TI뷿y^�<�J|�&N<P�JS�쳱�.D�
�`I�� # �@|�C�8̊��d�'����)TX�.	 g�9��q��sc �?������kሃ0�&*�Q�;�7�R�T`Ι3��ag�ׯ[Tױ��Α��-�C=�jW(�<��#t�'�% H�H-�l���#�P�����s�y�sQ#0�� ���:��x�� a��Pq@s�6��� �J��u�LݫB��>K�&�Ջ���}g~@�B�*���� 3f^��p�3�g�`^�WmF��hD;(�W
�+V,�c�������-��NU:UԿ������Y�^���O��1ǿ9�
W*�����F�f��0�ǹ;b��Թs熞�9����.�x����M� �DcqVᓊ��#ށ����)�@���E��.�qkW/_-�@�#BԚ٪VTH��DB�:��nq��,�S�(BA�t���PT��8�թ�t��2樂d�`�5]@���  �`&�ӏ���s6��hR�ahwΟ�g���&�у��}��[�?�R]xUH֠�O(����3߯)S�Y�M��F@xg����m$�J@���M�ڵ�ScG�t���k��wjs�z͞s�~�K�P��n��Nt�a�(�\}���d��#�a�c��Z�X���wp�S$����q�|r�q0���D(>;m[1����ua��;�Zda��*�e��4�8[N�ӏ͝;��ag�J�
�`��$麥LA��u���ӓlX�-gX�xKE`�-� /�W�w ��~��E�Q�ױz@�v�@¶'ՕԸ�w�������	g��ޭٷܨ^���������c�ЦMy����U.7�,*>�͜y��L9<DRT*���8i��H��p�@��RwG^������Ӧi�����Mw�W��V��s���a�&M>\)j:gɈM���٤�3�"E�Al64��.�|��7�u���8��q�`��7{�p�5Ny�k<�b�`Q����WųV�Ȱt:��.��7�[�n�xbsKc`��1WW�Ls�8��)D@.�B����u��Q�K:㒌��p�w�:�Շ��pC�\[4Ǻ+��&��j�^&�V9ߣٷ^��a��^���M:�Ѓ�l��:��K��7&�,��`��9+1G���4��3S��.x� ����z���RW;󮬹�]��3OQ�{���>}sѯ��}&��+����NRO1��!	_���͈�\a�q���\O��;v��������l��̆�̵��qDD���Ys<��,�h�kJD �zX�����V.j)t��ڹ���	��	������$����N���d������w�WBg��0O�	���3��.�|����k5��k��tj�y�ꃗ����F=��5��k��ѨR�Q)�Bh͌Y�4y2;�ĖOU4�W�17��C�8֫���7*����.��9fq�
�0��5TD�p��p�^�&Z��uX��q�'Em��c�]��>�~��,�=m����N����R�O���~���};�;`�y���qV����{�BZ�u[MB�w��0��'�Sr�!r��Mrh�N[7PL8�6����΂0��d�Z�`�J��ru]�u��������e=����_��^x�U�l��v���^�^9�;���/�����1i��L-���1N5�|l�O�����׋�.Z�ݖ������]�vQK���0��qN����������5�<p��W2l>0aq�m�����3��!��I����qi��vh��]�������Q�JS(>M�f̚��p�'��T+u���A�=q��n�\�Zu)��S��"��p��<�'iF�G�h�������l�LV�8�k�-�1=��Xc��xΈ��#���/0n?�f�p�'�.��@j������g��}�N���~�M�+m����<�6�ݬ*ŋ���ŋB�:�+Axي%!v�T(i�>y�L�q扪���֤��m֓O���_����J�:��C!����I����W��W��ߛT��oG@ئQ����\y��NL,�g��wo���+�u����X��'Z �>�@q�H��^f�NQ68 L��	q��y˽0it����=V�2��mVS�h-{�]g�y���f�������A��)+�)�*L���꓋ۛ�=F�q��/���;9�s=x���:��LĬ$vV8����w��^f���t𻁆�9�����r?��+m�6��?�q^L�P�=Z�4�\����̺�6G���g�jp��o�1�������Ƞͽ}_��>�{�c݋���0ǹ��e����scW��eID���.�4K��r�f��N54�U*d��쮍Kjo/�P��u!A#��͙�b���W��7_���gm<������ZY� cW̼��S�����+�9�U��|�Ec��'_��v_�jѨB�I1a�[8�zŝ��TK���|_���\fC��9�7��p|ߪz��vi�j�H�bSV�j^�BU+���K�/����*U3J��	�8W���5�����d��3�����d�i��'�A����,��!+&���kX����f��z�5�̽�Um���l��p��f}6�����m4�Ƌ���'&��^n69X}�/N����	䁺o3��������`��˱6�Y�f��a�bD�bY[�q����V�I�A�>�Mܖ�����#���bL�Au�4~L�.��]z�U�E�D�R��S}ݨ��y}]������f�&c�d,Jxq��3��qw�ׂv-��u��{o[�?��+vc�Hᜪ�	ׂp̸̰�[���9H�����ʃ�5h��vA ٢�c�~���Ժ5k(�r��r�z�*�S�ohQ)UV*]PEe�
�#�-���(��ʹ�K�<�'񍞔V�a� �����4�&����ӓ�L$��a�-j5׌ˏ��!k�~�y��<d0λ7��b�N�`�um�6�Ӷt����ك\�u���݋�˪���=��1+�6��5G�HUl��d��W;��3}����!O|�u1]��y�~�����k^di�Uk�(l��UL~�?��GWV-�hۨt�]�P;K�6n���{�Oz�v�c/e�.�N��t�Du�)�6���M��˹�������cR�������~@��y�Wu�Q/�H[���c�K[
�0�~A�6�n,>��b���U�xL��~haN�r����sO������IM���F�lV�RU��8�U@�"M����[� ��;k��h3��K�l��$�0Q)��>1	*�!A�	j(a7Ȉ8I�'��_(t�9 $��Z�����'� �qA���d�=U�l��b�]p�N��dbq0x�:��ɉ�Ǝ?ˀ�L~��K6��L{�;X�Z��j=�|Iq �+�^C��I�B;�XDlF�:�[& Km�h�F�i��XB&�.���m�t��yCO��g �\YA&X$y�ĭ"/�̟Y6ϖg��[�ߕ LQ��}�U�lST%^2!r�v��봹�K�:Y�l�r�d�qU*�{���	O��Z��s�x����rCͧ�߇2G��%[1h���]½���΂��
k üϷ����b��̭?&�C%�7[/�淿P��LU�Rw�l�ʤ���5&@�) <�d��a&7���%�� �~3��8��p���0)@��JR 79�8a|��\yw�1�9 ��K� �g�@1񩻊�)�xҖ_���xF�-���m���B �v�`��I��Oo[*Ϙ
ZLt�B�8��}�%�˽�~�\3��~�0� ����CF�G[��"O�I�*�����!��ܗPo��bĽ� M���:,X,T���; ̋E���vȀ?τk"K@��Bv$, /G}�4�+Ax��������J^jl�W�ܦ��M�$ �󅂪鴎<��e��ZM�.���WM5�.y�8d\ׂ�@�n{�����������= <��ˇ�9�Q�)&<��QadC��b����1� �؛��\�kS�j��?�C֭U�ܥ|E�[�M�ղe��kV����J �`���c�2Ø(v%� l�	 ;X�?�,3�aF|���9�&�yp<���
�	l  P� HS^�: nP@���H6��`��I�
�'���Yک���Ϲ ��u�v��~��<ٶy �̖{q-&�h3��Q�q�S�C�],, ��� <��*,<��s/��>Բ939�Ŏ�xN�'σg�,���^ 8l�c i�N_YHXmd�,���`[6�;���b��<{�gjA��^�M����c�}G�.JS�5����&�^T�浹s��~��z�[߭}�>T��U��3���9v�B��l���V���s{M��.B55��Z3���]f&Nx��+5�;O��φd�TgC&$k�����r���<B1(���*n��U:۴�X�G��"����L$۸��Ô��;?<��L�#�>w�)�U���ՓߨƦ������*��Z������Y��z0G�5�bM:�e2d�kA��2�`c�!�~� �l�]�:1��<��L~ؔ��Ӏ�1��<X[G��#�r<�@�8����y����� X�B#{���\� �xN��H�7���q.ㄾ��{����?m`���������S�9`gq��� +�8�|0K(�A.Ț�T�b���A���� �bd�����>g���g��u�xq��;��MH ?�ݶS�a!`Npm�X�I�,c��{7�\�bqp�mZߪ�v��}�l���ǩ���r�G�ι1ڼ9�je���VWwYM�Yu�t�:�����Q���Qf�|�]܋��X,s�`<ύC�)��e����������No�����4�|Otļy����/���ܴza}��̦Hs}5����P���Jp��q��OT�J��{6�L
ob���*��t�Վ������d@�v����������	�Þs�r�z��Z��S]t������^
;̚	���Fv�M� l0 &�6��H>��C��N�(X-�������W�@� ��f���0���G����C��^`ŨͰQ��8R���X8�@���� �˱�����xؓ�aV�7�����X!;=c �9�1ǀ H�1o�BΜ���&���ڮ%���{ ��XlXt�&�&�"�<Y� T�@�]a�L��&���dK�i}@saQ�"_�c¶g�"���ۆx��$ WՒ�/�-Rg[�Ǝ�j�͗�BX�t�ڻ�4n���v�mzmr��Z���U�b�++��w[6C��k��2 �w �,���f���LМ�#憝��a�&*�D�d��D���`G��J%��'|հ�0{��~���ζ��)�TQ��O1�W]CN�<�+%*��� ��#<Ջ��g�B7�5x۩��v�#`;U�jq��"�@�d��!?y�3n�~���j��M�[�:M'��`Vk�t�S�	��JՆ�w���5�� L�"|wu5;��	�2�=� A����dE^  �= fnL| &� 7&7�s`��x��+0cB0�`�� ���po�wHh�L��6/ �q�[�\a�,V�9���l_f�� Ф/����-Σ=��x�^��π0� g�q]Tz��
� ʹ�``�˸����3y.��p��EF�l����2d� [�s.L��3��3�9�;r䙳��o��bf*}�0h�:Ni��%z��_S�R���Ҝ9�駟�;�T����	=��K:d�������Ss�u�t(WGQ�d�O����5s5˷&l<�fc6���M��/�\kb��	��$yZ�&��e�}�	1G��r%��~��{����-�w_�baK���lu"@�R)+�n���'L�-�؀R�H�B�L�o��V{��v��F�� �J8�Sb�39 ہc/*�������)�Թy�����6o^���G���7d��S����_����JҖq(�% <� er�����Ң � Z��3Fd�V@��
�,lK�X�C^PX2e�H��°sO3E �g �ƦG� 610�l�@��!6Q �k���}��2 3�M�8�>9��`˽�D�%@� sM��Eơh��1���P��	�v���B;+���`��]@��J�3����"�2�9y�Ŏ6�Ok�Ȝ��\�5�d��	�̐?��5h� ���y^���?�+�l�KAx�KZ��UK�Jk��Ϳ\�{�z���ӟ�J�7��|OVW^s��8�DeӣT�H�2�T({03���GN��y�hO�ƳD�@V��ĵh<_�<�d��r��q<���D�geG'��:���W*�
Lx�A���n8d��Uǔ�Ǳ�Z!_
�,)��^h|��@M�vb�`GC�\<�a	�AD�a��n�4�z�:������78T�������N;P���f�m<n��ݺ������뀃���7�z���/�×~Lmm�p�Rզ^&|^ �lu
�}v~��&��ʢ�בpV�@�LP~�%�¶+d�JS�=�vu_�l��0��'��sڬ�c��)���ن�p��{  fl<&�:�~�xb0������ar�x�~ Q�f��G����1�Vo���N{i��/:|v�/�O{��H�s�#m������<g��$�����lwx�e�}�䲘�f�5�v����ыK�롅U,nV}]�����f�|�6ml�=wߧ�}�7�m�7�7ݮI�O�]=��R��d�Ą�{ĝv�i����(������a�4.>Ƹ����7� [s�Y�vf�c�@:x�g��&�q�K���{A��ٳgo)K@xb뺅�]m�3�\�	
y������+�q�����eU�����gM�`m04'��@C�`��j�đ�n���\F����g6��Y�A���C~%�|gE�n�E�?�+e�6����[O~��-[����a�{T��$LX͚u�&M:X�\W������=�j7�b�۔c�*�M0�����;	��������68��N�>������v73�Ë���+,3:O�x�q�l~�M��VK�����;'��teU���Y�q�9����30����m��2��W����Am �Z �Uf'����8b����8(�}6�N��6~w�`����#vx�c�˖�������o��	ҭ����N;I�m��9����T��{����M=�(�yerITQ�i�*j�02@���;�`*��8ϕ�Ȍ� ���������52��*�k��XC�q��@��,�D�`�w�5��s��t��a�Y㈫n:t�+d�[��A�!�uww��o�K���m����i���a(m�ST�Xږ��6ͣcѓ� � �O�l��7T9>�+_	v�3�8#�!��F������ǜ��+OG�    IDAT�+ ��ڭO}j���ԏ4i�x��wh����3O��%L���T�և*j��9��!�vN��.6G�m��N�X��@��6{d��r��"��;�œ��s�rA~�4l����s�����3�y&#���ʽ ,��g���|���Ά3�X��Ȃ����U_&�ߛM�U#{�9�?�JdO>�iƖ��N!�B�9����=�!��Ym�4r��zA�>������{YC�Y���SZ�b���Ejoۨ��Nͻ�]p�iڴa�>�/�_�ן�Ҳ����'t�qǆ"�
�d[#�Q�p�9��o���l�v�7�g��}.�5o��0v�����O�<L, ෾����*X���8��X���q�E8"�x���[���r&�}��9w��i�h�G�Z�`�JǱ�g�������t��S��w���Z&(����O���)�L�1���c�;�ٝY	��mo{[��~�{�9`G������������I�A�9��=�R��n�2�c��X�]v�>r�tuw�h��]p�uj�{[M�#f]lI$v�����Q�X�/��<t����'��fu� n���,/��|�sl*�y�A��s4��e�@����ф.d��	�1b0�������@;=�j�7�r���%���k�6��k��rl�����w�s����}N��5,��vm�#�ux�ŋ[��A:�%K^5���E�4�u�-�j�̓�M���_?�O��`�,��Oܦ�'��ik:$h�v�9���S5��1g:V�BB>>�<�����*����
��9�6f������9�@�߇gRL�e��t��;�뺩S�&����4m�L���������:{��Gu��}�;C��~��:;��
�xŬ�3 pf��`KF��>�h`��G��X_�@�%�53 �=�s-<�cV���chS�"���z�ձZ�<�kM:dM:l/��}�z������nVkkZ�*{�I���2:k�E�t(E�]E�]�� ���<�v>���F$�J ᪖�X����ʥ�V���C:�ijl��:�z��.=�41�j�}Qk[���L����جb>1���	���}����H,,���4l�̗���}�-� #�r���hD��W���	<6=،�Eڡh^^4@�4m|S�F'�(���J�J�\��;����
�؄'��]P��z<!j�i�6��N�!S������/�PHV�����%�ۅp<������?6�X��a' �����9�;Ǹ���5����إ����R�s����ܨr�S�GM�_�ިY��PwWV�j�7��f��v|��Z�gϬ��tF����.k��%z��QCz�T�М����oR]}^�tFݝK��W:�"�T�dT�P��v�b���0G`jt$��ؽ���`���7�	0��a��=*�^1{bv�s�5�X��и!�6E�u6h����������RK�l�����#�<rݎ�A�0 <�u͂����c��e�5�y�>��KTɕ�_��Ouw�H<��Vt�^fb���x1n�i�Y��P� gױ���TΪ��w�3���� #�4�#x��n˱3����nuu�V�ؖ�vR$k�U*JK�n�}�}]�6��	�>��532G`~�-�/T�1�����#Ǿ�0���/z����zM��%}����䓧�P���J���,��'�\Ɇ��L�M<��3qj�",�M{�ñ_�)�NҲ�Λ'{/��$�g��@�W��::�� q�|��l�	�����a&���OÄB���e�5o�m�s�1�w�Y	�c7�Z0��}<�ly����^�v�~�įU�%�/Q�a�?²��6A��*d����'}�8<�
v�����á�V'�Թ'������ Y�X��?�ca`Q�uVUPO~�~��k�3�UW�S6�l�Ġ��(�kR�C��I�U6�c;�R|;"x��@����;z��G$�+%`^��y-\�U�Mj۸I���'�|s���+956NдN�!�r%qВ�L)K�r�]3��π���K�%`i���Q4` ����7���XjL�\I�s�CS�l�4��\���8�,<�`|�;�	�'LX�\.�y�n�İ���+>y0��K=�I�8���u�Y�ӟ�{R/,Y6��� &:���!^]Tg� l������P; n:H��?:(������Fx\�$�jbo:�?Ɋ�.E=���*tC��J�;ܷГR:ۨR9�ԎH'�`�	;:"��� �����n���~WN��k�H`g$`~a�sZ�`�*��+$tmV�ԡ�F���PS���>5z|ؓ�2���$�48�z��8��sDQNl� N0�a�~�l'�v����û����\Nہ�>9d]:���o;|a���G`
\��.��A�j�C1��,�3��O+��<q͚���]Ӽ���'�E�z�;�ğ���V�8�L&�c_1�I�\���Kh���C�G��hv�qM �&ah�텈�`�#r�8�/��}�����"�=��p�t��?<�[{���,;T�kP�T�L�)ls��IBj�c.DG$�<Tt�P ;�<��ᶹbg&��9#ؕ�cn��e��N�K!���fحF��:��6�\M눩�(Wר�d߽�IB�P�$��[��Q�t�s��/��hѢ>��a^ޘ��8j₩�G@ؾ!;� r�����7�����IGP ��_Z�d���L�sn���7��M�g�w_�vas�sZ�H��ģ������Ǆ�e��T�0������E1�F�����>��!��f� 0�������#؏|�#�1�;�aV؎�f�i�P����@I�mՏ�oZ�f���;d����Z�d�2��O�	' |a(�CQ� �C8�2+�*�@LyWN��k�H`g$�5s˖�ᇿ�R�K�[�j｛�Ғ�w�[}C�
���<��������8V�=��	�h0G�Qi���cg��~O?��!��㏇�(�*k��8�YH�@(,�3;���9��	>0aGރ)�3�=��Ď�a�|���V������d�}���e�TQ������@xʁ�4s�=��Y=���}U�h(6a�ZbػR����Xe �L���0v!�;��L'�w5�Ky�)���i�Ɲ�e��1ʓ�̹q^TF+�6J�e2��K�K�����/��;�����*��E l��+��#������s^	��a�=�P��.ۭ+������ְMXH��ꐪSO���:5տN��(�kf�C�H�Z�`A o���>")�=d�X�D�M�x���;kҀ-�	�&�i!��%��q��tl
�0�����,�=��#jk߬2���.e�2߸��oVs�ԫ�?p��u���'x�Ͻ�碑.�0����~a.W�b���@��b�;��-dG*+a��=�	�� m�cUB(mm����Җ����%Y#횟}�R��Tvj���l�ޣT�Ki5���/��z��X	�V�	�9����\�{ߎ*j��)�0{�"�O��":��<�F��T�N��~5���=HF��e��B�j�G�M%͛w��>�uv�������+sZ��S��8U+cC��T��7"D-��>�����8I r�c@�;8�����N�ҹ�dġ����8���^1���3|��`@�&� �h.H!ף�z��.es�o�y���k� <f��Ec+�����!jg�}��;d=��ߪ��6��� �� �8V�^J��� ���@h�|�^P�9���w1j���"D����W��+ck\"*�#%,8�8��ؼR?����v�[�v�F�\�Z��[g��A�J�U�6&)�J' <�PeȘ�Q<c�ڀ�� a�;j}pL$���!x�}��#�-%08�Z�R_���*�ݡ���n�w�Σ�p����v���詧�뭚0� 廉��R�+��$Yc06�?~b��� + 's�'~v~,͊���7�9E�0����s�{z�?��ݗ�����	�v&&��`�����^?Tf
)'Y�;�nXA��5ƾ��|�	��LȘS?J�s���������z���a��}U�輙pl�v�\S����&8�!ܦ
۔O�&LX�� ��[�� �̜��Y`�0a�6�A8ؑTR.]��]�������f�#��
B�ٕ��>���T������i��I��5U	�4ү�����������Z�r�82A��#�	����/_JY�-Me͞�A͘�%�����|�a�ZӮ�o�SG���aB6��	c���K5 ���NlvJ��|���aV�h1?��o��0h�o��D��p{G��d�E�l�4a�9�{`��
6d�h�إ�z7	S;"��}���f_7u�Ø���ؽ}ݢ��'����F��رct�ߢ7|`��t���t�@���<w~c#ƏB� 1�%��x �f��}�C
�
��������?ݷ����4�v5���	��@�;���Oݡ�����ܻY_��{t��x�K������NtD�T��a��?t�z�����g�_Џ8�/�3���\t����xG bk�D�����t���K`0���׷���ݝ�R�-�߯3��6m�ܡy�>����/=������:h��*�K�P�.K텭���˂��5�*D�9~�m�з��H��Ox|�B�E�a�(�f��2�_�yET�\����a�r-k�f�0i���&RI�F�%[�Z���G��'��Z���~"L�8a�@���|ԡ:���	��+^�[��h��i>�����go�� 0�r��O�� $�>���"?8�"%� *@��j+�ج�.��,�RU��K��t��y�w;>�z೚z����3.V��S�ڒ�p�N3g\��SV6[��U*8�f��a(���vad�`r�~ ��ih���^Ԯt�.y�����70���Փ� ��Y}��o���U�ZJ�u�t�9����_�u�ݮ_����������?�9T�G���Nl�ٴ�����'l
��
iD*�O�_��onn�-���hB\a��m�Acv��_�4�'��wQ3��b��&,�u*~���e�ד�J]]��[o���iӦ��؄ǯ]M�Ɖ�	��a{�t�t����أ�Ӹq���p1�����?��`�&�a�AG1�s\�+k�1���3�LJYb��f�\�LV�/|�AE@�<Xo�Dz����(��on��j-_�gM�����7j���ֺu�:����z�e5�4��A�����c�)2��ׁ�6��4��]/���D_-�Woҍ�iD���F��|H����TԜy��Y�RG�f}�s���=�55�^�Ι�>$T#ĻB6]xU��}:0�ڍ>�1G=a���-���s�����:��#+�〯Am����C� ��]��%P���� s#đ�9�V>;�ӛ�Q����% <a��cʅ��ޜi�mη�yT��2U�7-��l����S8� V^�upN��f����F$k���7�G��T�{�VI��io�{1�ݖ�b�v�؄�֍��ݬ�z�N��מ��ԟV��SG{��j
�`�9+؄��\�u��N\�W�-R���"��1¶;8ݵ/���`y�H൓�� �l��zh�u�5fTJ��z�f�z�*�.��W�>���I���[u蔣�1M�1��d�^��0�
3�ܹsÜ_�j̀��������ĵ��i �d�;��8잏 ,ٿ /�؜	���L�0�g��qŕJ��9��[o�5Lx\�xb��
�d�D6�mN����1�����B�Pv�(�����xl2 0���#��@�]�B�	cv�m�qp��5�KF�6y`G��υ]<�쬑�1ݐ���_�{B���^G���:��m���s����؄{�VΜqn��H2�
�i+(��A�v�N�	�xG�D���+C���L#!j�4�Ϲ�PL�9-x�A廪7:�o�0�ՒVO��5�
��/��>��Ɩ�JSE��v��U%D-�Y�?f���p;s�p��͋`�
���?>�)��El� 7$�k��t��ǥ-}�XomD�wo���@8��>:w�܏�n�DG�ߴrQK��D�c�ʬZU�2�$[;1����!旕��sgX� \o(	Sv�84�������5RFWWO��^�u�{OOWXA�	'L;a���`�`�-w������Ru���K*�Z��6�;�*��4�PN+���sfhʔI��Q/�=�Q3�H��i*�8|��r/X�����Ȏ�F$��I�NHQY�V.	i�]my�4�u��W��oW:���fG������)��Q���Ja�V�$`�4����,X�Y�%m��k� 1��j���|M��/�7��p��zY�\�;��r��^����o��U�J���I5�;3�8�
��&Pώ����;4������ $�"na�ɞR�0��1���q�^޸B�\Y��V��W�I7h��n�}���^U�RU*KX]Uӧ�*���M���ԃ9���AB�9*����x�����H�l@y�5"��N�0�d����E��OiTSV^��t�a>aehl���T��Ln�R8�S9)ݓ��R��L�1�_ޜ��Wct��I�5�8�y�\�ak�6#�D%�b�͈��7YuXm|_��X�N�ӏ�~���+u����n�b�b�DG�Np��4�g�!W;��ǳw��ةeAqm����������?8��%������P��nP6EUa���F�Z�I�FOT�RV:���Q��;+=a4�8�@v�X�Y<�5�xa�ܯ�$���l	©���X�7*t��l����UU�Š92�w��u:餷j�}V�X�bU�$Ta�`g
"����-�y�0�dk4c��9�j��kƱ�����9��սE�|m�g۲ύ�V|=��L&��m��v�����k�*t�4Ä�ej�T�& 3e�h��r�7�c���ʎ-��8��1��Ât57/tX5SE)�YO?���=�P/���5�K���ZT�H%��Iv��sH[������PL�jmÎD��O~�`Ba��S�Qر�&(����#�m%08��li0!T�%5d�JU;���3� �f�l�0f�z�0�5�Tr|p�=sɅ����1�=c�͵ф�1H:2��ʿ�e��1q���s����L� �N��3����9�U;��M��|�'��}ͪE��0�#P'�
īIl����U��lA��@��<�=okU���!j0�r�]O=��
I��}�
9�ꛓ�wҝsd��8�����O+`LD^Yd��h�XW��f�#{��	��%˗�z�*���*aa�ʅ��Ad)�ޤ�R��@Ө�*���5%��{#h�	Ywwg�Y���f��&s	~$,�6_�q̌�ƌ>���p�&E�|��Zm>&�����;���W�)e���#���|��ի���X�A��qm���Z�N�	�(f۱m(�	W��ݪ����ڸ~�����rwO��+��P+�Q�J:ط���szm��Ʉ=` c��������Ӊ�F�v�,|�q�#��cF$0��&���p�C*vQĦS{���1Y�H��ԩ���1����G�=��W)5(��뫔X,���r98֞|2�Z�����kf��h3&i��c�5�Dc�#f��c��{̒{1m׀�k^Z�R�~�@�T5٢�/��f��+�k�c���%bVBǂ:���!(�f%�  �X�O�sN^]k5z�¾X��Ű��ŭ�m�_��U*��Jg�# <eʔ�6G�]��� Y���:f��w��,RC�p��	��e+_�׿�����7�NW^u����#�V�
Ŋƍ~��;	MjT*�$=�h<��|Ü�gBW�]'�I6>�1��6�������c��ٳA:h���0������y,���k�����Ͽ�Ug������W%pcP�����m�v� QO��X�<<v�&��M�`�<,?�-���J�.���~�(�_�\}�TNk�:w���`a    IDAT���G9�2I���ӧ' �#�����h?�7+��u
pf�%�G��q��w�z��N��A1�/�õ���0|W��Y���>�L�G.��ٙ�vN<v�����/y>���hVIs�\���y�r����FUK{hs[F�7�U(eB\=	��Y���5�xLHb�y%s=a�ۚ	�x{�qb�'� x��s�W~����&ĸ-q|�.aGG�*u��=氉'�l��|H�pt�qg��@v��$aN�p�Z�[���yW��5�2r��q�M%~o
Z˄����Ӫ���{�{���õ�����K+W�5}���jR��S�.'v9�ܙ�2irȶÑ��+MR��zW�����'C���svtt|�dlj��JaG��?�M�TiKIQ����n��ğ����{K_�)���[]��?�;�lyv5��kp�s�U�\|��������;�l���=nG�G������#�RW�f�]��[ޯ���%$cY����?��C&����N��:KeRɶ����Y��ɞn�i�1	ۙ>n��\�w��-��o�I���N�5�����keҙ�ϟ��2���5��d@�=�`K������x��44�w�"���3�p�2 �ٕ��X[��9�v����Z��Ԝ��iݚ?�sO�͟�Z��f=��Z�:�*ut7��\�t]6DI�7s��2E�
ay V@���ϔ���U]�>������|�eb�-R�L�d"ZM��[/r�N�-������F�����{0X��D�Ɇ��ҽ�1����}�xy ���緅�mӇ�a��`�����k8�$)+��|�2-Z�/��lӨ��n���{ީ*���G?����s��P�k>z��:�x��;�9�TnT]&�j%?(�������w��П�o;�I}���n���`���~o�mw_q�qSV�H�����τuk����0�R3a2� u$K$5|c;�iz���I��c�k�٫�s��wtv�Z�+N{�D�퍼l�
f��ک��\0Zw�y��9�h�^եw�~�z�-*T����<g��v�R�l0q*3�{Ad��3�-�[*��>��I�c hIo���m�3h��kGA�(�[��=F�w�~}�m �5���c���0�$S���{�!A8�pU����\m_���f�ܺ7����P18W�t�-\𠺻6ktKU���A���ܺQso����ȟ���[���iǩ��M�l&T%�M��Lp1�ZSA-�>>�d�� k?��$�^`̾��� ��cRi|�%�߻�ۮ�8a����q��Z&ӥ�M���۲WS|;�\/� ;�l��m=��' ^��p͆m��M���%��i�l,�t�N]m=����5a����懪m+W���PGw���z���^s��:[GN=J�䒌�
��w\��cOa�d�0ch���v�z:���Y�1���b��$}
��m���jp3��(ÔR���H���X�v���X�I�h�����HQ��=~{�E��ķ9H�v�r[�U���}���ѮQ�Ӻ��K5}��նi����&�ት:���u�e��ɓ�ΕU���r��j�8$��i7C���\r���;I��w�U����\�w̘Ì�EcsD6���=��s�a�6|�,�ݖc&L5@���\R��*���!�������pd�'*���+5x#(µ;#���|;WܞT�*�L����-�d˪��K�W����?Ձ�ї������?-�E�Fm�)U(:Bzr:2َ9�U��]ׅ��v�����`��̒Wt�P෽ ����''��&�W�����@̴������>��)���`~��]�Y�4i(�p,���� ��m�  �~�˖/��C]��4�Y�e�e:������������i��u�'g��#�R���i�V.���	T�2�؜8T;�s�:�#��c�F���Y&�h؄�Q�����xf0�S�{�����{�U�
�G^v�!�Z�,h��<��-a�N@8�K���[���!����aa�����l��ST&5�N� \���h�|^�öG�ap�a@!�`:�'e�舸T�A����wv���/WJ���+>r��Œ�����>���*����@u��}g���=^�<!4�`��5�9b�I�kn�[�q�$v�����@oi�P l�ؾ�a��Sj`�P�P���^����P6��Ȯ���؄��M@�H���՟\SJ)b�۽0DK�6�C�;��[����2GP[�[�\���657V4�+u�'+��~��g�������h��>v����T��Ov�	�l���0�0°�F��1�M�i͵�(f�: ��h�^��:��E0������7��7�����n�͙3��a-�~�U7�ۆ�{:�c��؄�J��l]F�[���Ïu:YU�0�Pi�0'������c����fwꩧ�z���8���/��{�e9��.�f�\��A�+�VL8SV�g��x�'�<y/u�!��˨�/k�ڂ���~�wfƣ�-�}�{���p�J=IȌm�M�!A2������w[�l���@x�I8�c���?`�j���qt�6����Ȃ��0���j�^-�m�{�/�dk��|3��(��o���n3~mӏ�@���y$�m�0����� z"��3�&�
;T,x��*���PԜ�.׌�*�+�����K��ǧ�h�����_�C4ԏR�@�U.�Sjm�1�����k�;���di�=䍲d����k��%a��l6���v�'�x��8�����${�Q�2�I?v�]s��퍦^��I�oZ�  �� �M� �����~�Lc�� �m*�6��@t��T�uvc����1w������c�=v��&�	so�f΀�%�\���U��Ù)J�M��{�Ǝ͉ݗq�Z�g�yI]x�:�R��T(R�>]o<����	�
��bZ}D��c��VL�wB�fǓ�f�m0�G0���1(hl��k~(��\�õj�G& 80VE��D�b�ۧ1���� ��18ԫv1��0��b^�z���_��ݪ�/��[.�y��b�S�,��ܢ��Ps�x
�r5��b��+µD��?�]�&��5YФ!��*8�\v҆�T�F4z��9��=�zꩾ�,��e���]
»mZ��9�y,NK�I�����3�l���z��a�"i���A�1x�#V����g��q�V/6�H���/���?�τ{�U	[ }�_[� ��N�@��1{7ͬ�w�*�jk_�Ɔ�TI
MW+9��x���o�ӓUUuJg�rw�6Y�nPkx�I�ϖW����n�֞X��)_
�℥;3)`xXM��JbL�H> �x�����g��6Ɩ��P&�>U�8��!V�X�ֲ��VD�1�}��'�%���,�Ύп��+~Nm�ĹB�կ
a�������F�]ñuu9
� �*�ej�x"��{�����I)��λ%� �O� �-�^��ܷ��\��I,ט�$~�$���t~0p��P��$���(̍�8���uu���~��}�qe�%K�����:���IS�0����j�(j���C�\����L�m�R*�jjjs��ȩ2N����\gW�g���ȁ0S�����TfK���Ȅ���P��Nv����ga'��  �`	c��M��p.�I��aA�e���q�]�L�:u�v[>��O��v̓�
��2�Q�(�?z�({�њv��Z�z�V�\h���=z�Z�^i���st�ݖ]�΃��`�l�	�bOfu��y��a~FV��7�����s�;6wl�eu���O��Z�v�Te�����ƌ�C�ֵ�R�*+5�Q=��{ϰ��{���ޤ���'O�؞h[ؾ��l)~@mY�aI:vb�J��!^�.I��e�"���8&nG�����&��+�)t�A�� �j�'wr�d`�a=\{7:L�c;�(��bU
q���`�b��$B���6�j�� Ό3#c��MS��'��"c�&�<b�N�p뢄����2�<qó`!������_�O|��8����6?,5f�-q���/*p/z�L�Ֆ
_�s��U��������=�+��6��o?�Xجa�(�D�ӄ��e���w��ή���Mx�Nz��zݞ�W&S�8��qT,�o	�����K�ro^0Q�a����wt����;� ��Ny�P"ֹ	���Ш�M ��/��!��x1��&X��6��'�%!ʢ��� ¹�G���k��'�]�`K�+0a�C���#���w���`����/���\~X `��:�4���J������}��U��a2�m��0-Pi��b���_���m��<�`Vm �-�R*t�d��*;C y]]�@����=U��/{�'gUvf�i[S6��:1�CH!�PU:�ˇ�AA �PE�E��B	5�Jo"Z�	���u�;��y�ݛ1����_���o7�3o����<�Γ\�e�!1	����Xc���J\�?���V��/�9�M�;G߳EwY)̼6�n�1�YW��ݯ�Ɯ'����8Oĉx�|l���1�
�LB��.��m
����A�o9��Ka�M-�7ӓ�GI�1aס���\���}�SW`��-"��.ס�Y]�J�	Yݫ|\��/.\ǒ�e�� $�]�u%qL�����qt��Ɉ;6@Ι����(�����g���Y�q���f�v������"�#�qEr�������ΊAXI	*r.����f���?s�!, �8�	�-�;�WX�p��o��Ƶ��Vj�7g�IsĀ�"8�����s�_~���٧���H���xI�^x��;��Q��Ր�9�9�?��!+��G�l�3*�E&f�E?��n�����OħL�p�p���[R��Ƅ���1��n�0l��x��iX0!2�\����ׁF��������:o���τe������K�������O-��|4��b��G�i�#� �͍`��)�x�|���4�2���cv��B�"K�@�A�<�aw���d�b�n��i�W(tXk���K;��%׽�Mhg��bN���9q1;���'&�	Xp�l���Ĵ���F��3y�v�r�#7Q��h����u�����x~�)����-��Il��t���p��Y�]���������M\~^��B!�O���g��j^��KznceׇRU<�����a5:�qH<����:	ܦ"�s�p�A`/vk��W��6k1o��;�2�x%A�[�S	�k������\_�by#����o!,��@R�Ϛ���	ekκ/��B�4��phqR��&K=�s��:�����&��_��5�y�d�Č]w�Ç7}VSY	���6,�B5���O�In�$���)S���^��)(�㱻ϟ8�Ǜm���e����[q���o�gќ[	�4��p5���H���^y�v5..�^����T�����e��鲛�c�=��6����(�����o��Ád9�	d�t�qqˣ�����R焍!��k����s�Q���B.��H��#W4d���>Y<G`󻓁v��0���um��i�S�Dt���a�d��N�E&78����Kf#UE�t��X
�{oQw00N)96L6K0��"�O�}3V�\�@�G)��~o9�c��e����<��F������T�0�D��ɘe��N������ۏ6�U�Ϧ❖Y��j�MQ�3�Pf���-�)�h�ùm�<�4U޳���˷��E��7�>�6T�"!�yw�&��O@��κ�g�I�):s��Yleˍ�)���E�`�M±�~�3am���ֱ���e	
�����,(ֆ\˳|�`�e��6Dm-�J�_Ѱ�b�b�$f�6LwL�i��~�3�u�Lc$�<���������_}�J�e�,�����7�4���0ٽF��׿�9�;��8��2�}Sfu��0��X�΋.��na����?����	��m[(9�{�9�s����"2!	�LI��JiBp7�JoaýѣG[�w�)�y�lxI� 566b�ԩ֝�裏ƨQ�p�W�.��ó��egJ�)?X���t��{�>�+�Φm�p��Yh��G��6cCe�![��P^�![be�N�pq�j Д�C��T�0�����C)ӈ�P(f�;{����,Í�kC $��������9b^�!$�Vf<��-����6c<C.H���]��.����\�%Ky��(����N��� eN��D�{<F�Dc�H;�sa���%���P@2�p�8S�MvW���L�������ܡQ4gn�����댚�Mn��p�?O&�+�ȟ��ʲ�9�'.ŀ�Y^?磫0��g�(_3�Y�,��ٹ2�Kõ�2�J�S�'����2i�*Y�Ry8IT"�d�o��ZfcXB,pL���'l}�Q��䇡��m��E,p#d����#95c�2�aS���8����ǒ���޸֙��O���� �,�ʉWd�>� ���_1bw\x��?�V�d�Esn#s�qm3|+|���������3?C�fe�Ձ�d�2�������"���3L�rPi^h�A�t�;�hM29�P���n�B���k�ΐF(���@g>v�<� \D<Z�[��B&�;�4f$@L��bY�$�vg���AT�[��}����t�71�yPd%0ǂ�1�x<06l�/:�� ��W�dO%�l�fs�NB1���f+e\�u;�N�عr�	XB.OO�[5�B�͓��e8qL�\+E˱�%45-� ��<i��5�g���NOfb�����j	dy�sx9&�{w&���
��W�{�F�nFZ�Ӳy�/c�9nv�n��5\:N��-��*��(9& Vŭ�T���?�.L�t:�{~����@'5e��x����:	�1B��M~_,��9G&����|5�<��:�1:ta��� �5(;�wY}���y}��f��,T"�CaB� S����'߷�%����*������q�Ɋ	��gZ��{y=�2���;v�������UЋ��t�I.�L!ي��嗝�X,�h�x��d���z�ͭ��X�.8��n�MN8s��f�V�n��9�6#�a����}�*(��wN�{��9�xѼ!���mg�曩|�4/��n��L -b~�i-�4��N8�{Ԇɐ�ߘ����tP�RϪe������3���O���մߢ9K�vʠ]r�h"�tXz�	:�r}�R������ �@eig�9&�r#��z�������O=b�$R�u�IUaIK��/�ʹl���mns s��4��A%9�ts��qV��%��>������ NĀ>=�@o��M�,Xf�6O+�w�f4�B��%�h��ȤsH�T[��6��Ǥ�Ǆ����K`�����-���X���bsk�ѷ_O��vC�݆C�*E�cP�ˆ�����ظ�D-r�<�j�1|Ӎ�e;�ܷ6�"�!�Gj0o^#>��3����������ݕv<òsѴ�(����·hk�!��6��Z{�(�l�"R��p��7��#H��fb�%��Pz0�76�p]�76�q���Yb�N�)��%����ȜĜیJ�x��У.�|��E��QJE�:�Ut��;g!>����q��O?9���4�ݳ\:��X+��ǐ);;��<�2ea�h<���� 5t�1D����&�u#�Aa�}Y̼:�H����B͗�9s(����H�د�l�N=��M]n��E����N��K~����9�x����;����"
� 2��s�>�[3�X;��ܹ���۷�>�n�b�Q;bܸ]��?^���s�	r�#�!P0v�7����Hy����,й���h��sg�Ճ�Nu�q���������>��c���ꪫ�5�嬑�T9�:��	Z4��	�?*8��꾻�d���i�jg�0S,�A"�g� g��x�5�$c�C47��F��d�+�УgZZr�b����_`��2�L ��{���N�.z��Ҵ��uJ�(|%�d�s5ҙ���V���_,���ev�5�<�$\�\1m��	^������e�����p%��    IDAT���"_�p���}p�٧b�&k"�ʡ� �L��Eʱ�b;jkz�����^�ioʹ��h<�w ;t�egS4�B���w��Ƣ���-x���n��6���@�^Q��D�Һ؜dEz�I��)�t�U���o{��L�Q��Uᢋ�ða�!�����i��"��"JQ�o'0{V+~��3��L]��^=�8��ð��۠��N>��_o�����Ǒ�U�W߄�S���O�9zc�q�ѧ���:���ɍ,�i��X���p�ݏ��߄L��G5���ß��}z�O�!�.搨�E&]v�E��T���᷿�f�Z���1c�G������kY��B9ϹYlPfr�	���^\���ٯM�M:�	´�����YSr�If�8��~{�,Ʉ�|�}�w:�h�I<���>��S�a�� Y����$#vQ�B"�|�9����v�'|����]4kR��y[�4�6�h8=����VA� �L՘i,t��yʓ*p$�e���	~���,(A�7��gJ�
���79�ػ馛:�׃�j~�Xa�:\���,Y��c��V%GÜ�T��gc��F��i�(z�^��۸&�b���j�z�q~�r*f�`A}���8��q⏾�d"�0��L	DB:G��������<Co�5��q�Uȴ-���7�o.;U�EDb$�=Ē`B�:��96���}�M�?�*,\�A�cР^��տ�F@UMK��B���%KZ,?�mB}�����y8�?�g� dM�h�?�;�\#�|����ȤCT��@1�As[�9G�~q�p��Amu�\6�r\���У��E��I�si�riԲWU)@6E����wN�E���b�^�S�������2��t���׺���6Ī��a��-8���֜4pC���y;b,��<��zd3�9]]M��B���5ho���s���}ɮ�6ဃ��ŗ�eV_U5=��҄H����$r�fD#Z�C���_q��? �gDK	��xn��r4� 
�PU� �#yh!�E�Q|2}~���a�Bnp���5�G��/\גDW ����1˰N�3�W�R�+�>�� y�G��Z%0r��QG6K�!A�~+̑�F�ʸ~�Ƈ~ءo���������=�S��;�c�Qq�a��*�-V]*���x|�ĉҭr�	�i�?�:�2B�䌎���:s��?�~�4a: x1��#;�7$�P�T�p8J���@�T��M�j���hq't!1α��\Dw8e�H?s������y1a1hm"b�_�u�)�����z�U#�m�5� ��C*�ܹ�0����޻�n=�[�a�u��̚��u���q�DZZf���cL��.�0�����O����ת�&Ç U�B6��g]�{��+°10z�!��Wg�GC�X���2M��1x���zۍЧo�m%<�ī8�UXҔC6���5{�ګ'bذ5-�z�&L�`f�^�D�
#Gm���kP,�ha��#|:�yV�����ӱ�ޛ��g�t�^|�~2˼�[l5n<��J/'�����Ȁ�m�&���r�� �x}0�0mm-Xc���醨�AP���;����X���q���a�-7B2Z�3fᓏga����Mb�m6Š����=�Y_���C��9!�R=�f��3�����BUUm�Ux���1�3����o���,"h�9g_��S���,��"|{�m���~�T��%L�����4�J	����t�:����}n�4��t��Ym�h����5�ć=���\�Ӧ���K��l3bK����|	�ޞ�SN9��f�h�p=$P��A��Hi�_g������qq�+.~%I�좋.2y��k�5ف�ε��q��g[� �F�>]I���d/2W9��Lc&�Z��������˟~b}�+�P�Z.�b�;'N�����?cH��_L�ɶo�L���܆�=�b�}��A��5.V��r�)���r @48�*��;$w$F;P��K��?C�7��.���p��Q�9?TG;��&�AO'�"�4�d�c1��d$��`.ǃ@8Z
Odp͟.�v#6A.�Ƶ�\�{�z�L�d�l�)�8�x^k >�t6�9�44-�6}-6���N��(~�Y��������-ns�o5��c��^���b�s~~��o�ek�JF��f�����ƚ���������Ghoˡ�z���18���Чa �|�e��G5hM�bР:\s��>|]�����<���hivyc����~�t:�c�>�L_�b���
??�T|��/���)�������K����V������{����������)�DX�>������Ä��_y#^}�V�y͵{c��vŉ'� I�r��8�j�Zcu=�����м�	����x�����j����Gs ��>��Gu*�|�A2Q�T<�?;2֢C�L~7�x7/\dRĺ�Ʃ���ѣ�`�b����	���=���~솸�Hā�>�<~w�x��/�0x@_��q�w�������I��o�F{:@�*�~��4�2�ѯ�f.���G<�̋h��|���Gu �Yo}����ޯ�����t�0�v��#1�n`	K^U/�}#q�V��KVvmq�Rz�߇�0�F��ɻ����DKZ�*�Đ!j<%	&������E-�Y�_�!�.C����'̰XFr1Ȁ�r�H�D���O�֌9���1��ɶ���,̇�S��2�v�c����{���a]���29� xC���!�exژ1c�ǝ�;o������3��Fq��%�s�YҒ�뮻����4Ox<�QҲ+͉;�9��K�Y��zEX�M����&g�:�z�1��`ܸ���k���������j�`޼�h�_��O9�}0�,n����%qsƤ��8��#�����s֯���o�&5������������~���/���Q��ZD#E��.~q�9�7�?.��j\����,�b��=
�����1��٧_'��$�-d���^����0|�zx������}�a1�"Wh�O�8�]c/?������tR�)E��s~�������<s�8ӢX�aqS|o~y�D��q�����?c�� V�&��[�E���e�^�{�~
�4��#�������?���C6ğ�<��ş�̉T]\�s0f�V����qٯ�-K���ޞF���<O��T~���p�yԉX8?�T�^�6�}�I8��=1�Ïq�����g��"��2��k��췿A�Ǚ?�S�>n�z��{l�_]:��/�◗�_0�)�$��x�6��.9l8�L�Ɵ�G�"5���֐�x��̂����p��+P�Ҫ`�q5=����}�݌����s0oN����lQ ԃɄ�E L��ײOθ�y��5��Ck��K/�O<a��.�đb
�$��R�rY����$1��u��� _r�wՖ �&>������z�vN�XG"�0��5q��S��7���k��7������t�Tס�.�_���k�=��:k�i���O]3���y�^Pi�t:q"����d�,ʜ ��3��w5������w_LFN0YCF�������{Ȝ<���X�I�U؂6�Jv&O�d���:�Pl��ڶ�����>���o��C�����h�^W^�'��һ����p�i��\��	S�~�s���`�� ل���;`7�g�~��r/Z��[�������x*�)S��鍨��l�� �G�� �=�������	�͘c�o��:��ʘ��t<����=�V,�U�؊ۭ�]v��By����x��O��=�z���N�ƛ����x�Ǒ�31$Rq̟7]��{wD�$}�9�v�ݦ�&SQ��iss�V���;�'����/2�Y�Яvt�>Xc�@���?pß���y�{��:}q�O�ƀ�x����g_B6�7Y��nɒ�a�15f4��<~y�o���_���Jओ����73g�#�����
�B(�h�B}�*���H$���C��ǟ2���6�}���/r�y�������OQW�a��l��y��X���6�c��������@x���8�'G0���0��� R� �@u7�F��ƌ���M�﫮�'�q9s�1���%��rK��rDe�D��EI %�u
�ZS$I���A�c+�%�����Ep$8��O��"�����~%FWP�,*��H��K�@[�K���~֡!�f�C�|�U$)�b��.���w;�?���\�H:�k�^���*K[�e��H�e0{�\�1�/e�H㵐�04�L���ed����l:?�L�p��Z���~�;�ŸH���5N3�������mI!+zМ.��K,D2JW�+&,JfN' �0Lۍ���ią�[ٌ��̌�\��<둘�a���;�Xlfu*�	'����ej.j-�!��X*ЊR��
�B�5ep�ͷڦ�H�=��[l����e�!��^��
%;�'�mv����cūo��X#Fl�q;�E]}5r�64�����X�Z8Ya�#H0�-���>�*��y�;dm~�Av_�7$��%�d,i�0�!�K�����0��|�-6Gz���~��dN��C1����JAU��Rֱ�\S�����c���a�=v��^
]]�\9�9�k�g��h�T5�z�I<��S(3Xw�5q���G]��7�7��_�A��L������,bL����%QW_�}���bNU�&)�N��u��IV�"��a��&���x���P]�n{C�1p��I�NQ�Gl���N�P�#_hCMm�eT>�̳x�o/x�i��ɣ���י�]}Wk_����(aE������H�3}G5UH���nSK4��G �c�ǣ��r��7�҄�Yeg2i��(7^j�����r�A)�H�}�9���[C�Ȅ�͙�F���ie3y$Kq˲bg��F��vێ�@tj'�%\��+Y�?�+Qb:!���ܝ�\`.vҥi���;��LX���|i���o?|�;߱z�<�@W�&���,'�o��{����|&�0M�]v�	#G���{�P���
�X���1�ic��.7�x�̥���ȣG�:��T;0M���Q���j-0v3Ӟş�x5�45�Yz�!�c�M6�D�D��ô�(�j{{K$��G�0�H�}�Nśo�D��a����hooEmM�|ȸk�YSRr������g�J��Ͼ���z޲��[-x-�r�������L�̤a�X�u�]k}�^=�C�ydŁ�ģU���N�!��1��af.d�����m�[>z�Hs~Qv1'pZ1�L���X2�x�������G�X$e���\3jj"V2'u�z��Z�03���]�[n�dCF�q�!Xk��(�]-�|ԅp�r!Xl(ɢ6��A[&�|���w��=��M7�L���8b�h�)茲�����H%��w�Y�)NX��-����kM-;��s���Zת)�26]���|�2�8~�R�E�$W�B�N}�׵�n%g���H�k��GC����s���;�k�3,�8Gi��^��p2����/>�[���c��Q*o��jy�ąQۍ��oiT��7u]� oȘF�d���E�I��aLa&x���f�>c��-�,���O3qȄ��T����yv�[�ʿWFX���06��λ����0[��w3�ъM�ooO{��2��wϾ8�cгW5r��9IYt�]��ɞdɽ�T��I����Cs���r46�d�����43��h9���&�4���g�ex����B�؆v�	;�ݫ��ێR��[X�n��W���W_�#�<jbk���q�Mb�vc�>�V�%��/:��y�����OV�&!%*��&A��2� ��;�[/&��z��������0v�]Q
�`� 7�(#,��Ӳ�-6�.���yx
�b묵6�8�H�V��4�H�<��}۞�Uch��'0g�b�1�n�e0D�����A�LCfZo�Y�ш���x�Ld`z4"hko�=�M����7��cϽ��[wT^3�>t���8w�RLRJ �i���?�g�}��	slx��#{f_�W���E�$�I�fh]�؈Պ\�s[�1���,�L�Y�$�>�E��A-�?q��@,�:��tApϹ���ne�C�?k�~?�T�ό^[�b,���ײ�gRv��0U<F ��M3Ώ�I�X�U;b%S��)b�0�$�i���IK�`� ���d�(myUO�/s|MM&��Qc��.��B����VኺS�'x�nU>x��0�d����w,�{�P�f��M��S�*���b,�l:���x5��̷B���{6�h0ق)��x3��ƺ\�6,PJ���x�W�۱�.���ݝ? ��5W��^JaWq�����w���GQ,�0x�z��P]Ͱ%��:pP��Jt^:	f�������Q��Q�C=ܬ)�"��X�,�+�t�v�w�]6�8�;�;v�
�@b��<�Fj��]�&^<��sx���a���z8p�Cѳ��B��`	",�hŜ�BM����1k�BL���z$r�Vt��/�"P���]��8u�b`R����<tޚ�������`�-G�gى,q�R�yj��t�C5)�z�	<�<#���)��V7��>h+���X�"C|8J�
  VY�hԞ�"0��S�	��Ĭ}�/�*�Q%r.�2�a�_B�y��R3!3�M2z��/��Ej��E���w1dW�fk����!���x�*�n��\Ԅ�g�6���;Ժr| �������k2'@ǈ#��.;u�׸�0k����\55�V;���>�t&�k�ջh����j���!�Rk��z�e�o�|7�)��X��s�!��Łi�g����E�$&e��5&����:�_�p \(�1v���N�:�-���5�\Y���_���NE.ߊ!��G�J]�BV�rV�c���X91~������N�Z� ��p��n�~J�r��e��E1���]�h)��v�;�0�
Њ0RD�M�D ,3EV���A{�ox��Q���zb�}@C��(�Pv ��v��Jr,�4{�|�1�.4��X����׊�S��2�T�t�rW���@ A�<x7�}w�""�b��lC+�K]�9S���u�ؼe�&"x����⋯�>z�,%s�r��^��u�g-'<׺�[��t�D�H)���"�:�i�������*0}]����~W�2Y�d¿��/~ԭrİ��f��ٓ��i2�@�@���m��紜�dҨ����	\��:�/O���f#���Xd{d����T�e�����oO8�L�%���"";ﴃ��O�r�٬�?�0�'�|��������'N:�x$R���E2�@&�C"Ve��`,w���D�=�o��g�GU���{ ��a)�"� �O�"�Z��=�-�*�?��|�D�El��6�c�q��zư�Te0�����xO<�(ҙfl��z����0�.�qԚ�������Ł�o�h֝���_�>���՚����u�ݹr�1L�4	���9'�����a���23�1�HH	B ��� %��ګx�ѧ,Ds���Ł��L� �M���+0�w�:{�,�:�6��6��G=�w?c`ٴ�$�"f�k5����x�-���{��p��6nl���	+��Jo&aD	�L�ȣTt�V9FO}��K&���bC���~��0֊�$U"\>;����h����ҤŬ�m����9߉1���o�r�y��K.���
~�g�{-�q�@�J�\� a %k�����H%hT�?`�@�Kf��KS������J��C�J�_��<Mؿ7j�����:��KC
������P��*�;�}�|���"��{��O�z,2�8k�DV�>�:چ%.>�����rf�j4)�a~Æu:)��Z�h	�@I�d�-�G{o���Uy1jv�aL�ȶ��:�߲�G]8���7^�3�<��v��z���}͂".]�[k�d�%���0=�}Ѣ���Y���F�:�k1E��[LK3"��P.IF]\��    IDATO�ܴi�%���{�յ(���61i���0.�*av���x���:���?�PTW�L
	�1�y�e.l"����3q뤛��i�1��?C�Ym-��y��PaW��Pb='�����R[U2eN�-�����:qƨc�ni���qh9�C�ԩ���^� a����X��^_���V������'>P�v�S$7?��O��O:�W8��|g�_U��Ap�������[�"+�Za��3&��c�Ǆ�@�L;�����r}g��8�J�
�����:��v$�I+9��c���ϛL���X;c�]�2	���+��և�&�5It����~�L��\CC_k�Ds�Be�.vR���R�|��b�	sF�>�N|1s�1�C:n���0z�XP���ddtƱ6��g����cx���p�[c�]wq H3Z=�:c��;�i�/��"�y�)��6a�����|wo����i�ńs�E	�w:��;&̤��o���fs��0x�Z��v́��`�\j�cA����`�;����v��Q��F�n�:�:4����x�W_S~�tu�Ї|� �ץ�%#N����Ps�����?~��{�/h�Ƞ���m���R��G�U�c�>Kf��1&v�=���!��[��-�ڼ����\��I,��4~
"�pK�>�����_�waiƄ��L�(�b�7 ���^O�����F��'�`�����U�
��b�>�乕����?��n�ދg2Dm c@��� l�˝'*w
޴
t�������BVV�~
�gU�A������u�T���d��׹x"Țcs��#)����@`�<g��aޙ��y띗��o�vۍDM�7�"�;��,یBgqmV$���v����|��6����0�5��$���='im�K$�� |{�[���f���κ�p����$A&�Yh�����:l�����&��ʭe�/F-8J� ��:�!�����|�m�PS�[l6���6p)WsN��~o;Ν�ޙf��'�����:��b���(Wi��R���@&��O>6g(+�54�[lf�4	�iv��|�"�ո���z���4�୷�FS���l�a�ӷ�1ב$�u]Fl�c�W��ioǻ��f��߃�\Á|YEp]��Ȯ�5#n����������ˌ�܃0�,"ʝ}	����}��+�o��6�Ë"�b�>�7������w���>+�\j��	&�ԭ �ى?ԫq��u��1%{���s-�����v���)Mƿ�=Q�j}^Y2~ڡ��ΤA��͔�8�?9:ƃ1�1.�"�S���5��+6�����bE}���L�B�ь�l�����v��&:�Lg�p(&-�>`�VTUV>,A�=SDUu�����QưMҊ)����k[ښ]�*5���3M\' 깱:�cîȓ
�3^����<��	�S�����0��=,�M)�oG,H!
6��Xl����խ���uD��@�E6�⅝%��*�=�v�p��+shl��64�%Y�k�i�a�."t�#y�-WQ~?�X��Y��=;�7Yk4��k�8vڣ����
�	�s9�9�)WX)� mmtF�.��"C�z���;V���Qu��#X�Y������8��J�}�O�ӷ�eY����O������ar6g+��D��Uµ�V
Fu�7����\{#G�+���+e���H��i��X��~�Y	��_���vl�C
�r^}�cuG����r�t�q�c��/��u�y��Gz���g:�4K;j��v�0����`�|�g�H	7�.j�	�e'�R���s���˭(���R��Ҟ;�
�w� P�K�"��pz�����d�K�#W��%���ʛC��7�-US�w1͝��ܚ�l�c[���p|e�	��u-]�}W1��h����z�����]!a
Q(r�3�2��QZ��}�\y߹���y�h4���	N�V&LM��a�X�av��!@��I#S]z�;k,}}�����^Y dE���Ү��U�B,��n�:�@��emB�{>�𿿬��i���X6w�������0�<�\|J���;�ry�]�.!�+3_*�ϲ�>�,Ӻ������蚻����o�g��i��@�oS}~��|�h���g�>��j|�N��RZ���τ�ͼ���:zy L�/\� �O>1_]���R�v�m���[�B�&O,�ں���\+�,|���	��]�ݲ��r2��}���X�;�騩�'��D�s��%�2��د��WW����_����9���|�>�?s��k<T���-P�wĈ�ch��y%�O�c���W�|�&|�y�حs��3o���6���4�r�����)��O o� ���=|�lK��nQ-�~�&�׽��YWLjy��
<W����8�;�oو�빗'��^�2?�u���l(��X�s�Y[%t5?���|C�,�T9����D�#T�M�$�h�?ʟG�/!�X�Y�ڴ?g���R��{�'u+3m��B�	��Z�</��k+5-$1�J�݊��R��`�;�����}C���et$��e��������|Y������q}r�U�Sy���돕�/�[lV?�?��_��+��O�8珈���	l�3�������
9��F��KN��R�,��s��I��֑�a�i%�w�7������.e�q��ޮ�F��Q�
C|����Vf��_���W�����W͕��(��sU]���"��b~0�@T���7���z��������r���խ��g�v�X��q��ܭ=�6��C�/�u{}�u��@�2�XN�P0�d`0�LqxLd��L�L�����Ϝ+M3��W5�W�����Y޽�*��e�mE��U�~oY�te����o�g�.��{�:��M�n�cޏb��STWm��L�+�%�7Wa�:)�H�2���,@ƚ�Y#|Sނ/i�|�b�H&|�E��[Ax��g�װ�Iu��m±�Ӏ���5�ʾ1/~��@i��a�(�]�|��T9〱�o�5e9pl����dG���T0^ނ�	�������u�/ouu��:��]]��t�	��*k��ݿ�wI�Xs�䎅���&��}֩a3O&�̤�^ͻxh?�B�	��|d!%f/�>_�G&P3��UӘ2�^s<��=զ�@x�E]��n�MN8s���f�R�k�jQq��V ��1�����f�a���V{�`�!��y&o�i��Q����,+Ț�
#Q;i�]u��]�۳Xw%V�g7��.��O�0������*�no�����#�F@&?;�����	�lgĵOF��cc�I��8C�&�BE�+,�E�`�`�5��B���bb�AbI<#N�K<�=U�����y ~�\�-�ܲ��<�֎��S7�;o�M=�V�PB*�B1��v�l�]w�Śpr� �U�y�BJxAܱH�Y��Ay��g��B��~rg#��L�gђ�>��w��3����*w)$�������J㑘��v�4��`����X=�� ��{��h�����@J�5u�T�u�YV�N���׋��'���'�"�Na{5Ue�3�?y�-{b� �?Or�k�q��*D��)&L�^v�i�4̟w#��D��
1�1z��ǖ�l�-�9VJY�m?|�]�D.��7�Ϋ�9�2�Ѹ�H�э�{�<�䯹�c���ؓ��m���G�?��J�p�k�M�_;uV�m�����-��.��<�1b�=����=(Y���+�4FK"'�� I�H�j����*J����ĺ�C��J��CI���5�᷑H$O>���O�V&��N:�i������0g=��F��9���z�V�a�м�	o����=�
��0�P?��7�B*d���s��hj3ou����47�ݔ�̎�,���&8���oM���P������zV���~H�Ȅ�;�<�)S���W^1��l�w4)����aGr��[}�X�/�j��v����e�[�8�7��|Q$�$�dƊ.� �A�}���� �gќ��m��Yky�]����i�ѧ���[vA*7I�+�W��5��;1ی����R5xj��A:��#�	Ҫ%L遍?�P�;�\~�pw�����3���#��� ʾ��%�p���Q�$��_�����2�
/��0t�P+JФ�K�!�v�������}=e�w(cЂg�]2r�����ly����� ܻq��#�m�b��Sb������Ǉ��?��#��7�~����y�d�܁�w�d���Ȇ))(�[�+�Ѥ'��l�i��&[%qP���Saq|�����X=��#�g���;�Зv�n�ă���o�%���('���M�GL혟q�Y�
;#vH��(W(m��S^��x6y�d�)|
�0���<��s���[/�2��Bǜi�o�/�o�Z��B	}k�X�چ<�ק�7w+^$���YQyi,�$��N�⋀��3�4�=��y;��q �w+��������d�qJ�)��|��� w���ek�gW����׎ q�k}�]v1ٓ��H���I��7#���0?O�ψ�A��Ad�����^)��O,cH-ϧ�3C�Ȉ� ��N�9A8�M�����#F,�2��%�il�!Ѷh/���N����/��q��oܕ(^��r�� i��	e��)�[�k#G�4`e0��;��q�g1}o<�!��t�I־��=w8�<�����`��Ϫߙ��Y6rU�q�qW���pHA=�@K�E�� ��{v��������"��ȓ-��s��̗���@�Cď�%&n����o�u���������ގ���b�L��s�9��
��ƃ�̽!ֲp;�`���c�=�������g��5O���]���y3r�|. �勃�}�-l� {�-����;������8h4'�B����կ~�O?��cpy����ᦩ�����.���R��Z�l�cA��ˮ30�Ė���x�ڳ�;5�/6h\�� �M���u�*��+CBW6qey��5O���^{YtgX+Ca�W���β�ӧ���B�����a�S��B+�@���
'�J��$~�	�%q��=d��AxqӒr��A4r���N�V9�q���ϻ�>�ގ!jl�2b�m��|���2>���fk����x#�q��͟8��f���r���;:2�)����8�ṣ��[����}_q��q����zt���0�l��;&��^w�H�QvSP1qW�[�r�B��Y/�Q �=%��`�)�篁/7�2�_��LE��s]o��&8ꨣ��&����QF�����]E��u�]�鐣����'Ű5ʜ���v��9AX	�Hi}�w&�͙7���,����Ϛx�O�n9���5�1קq&�5F�!��n��6�g���ן3&LM�J\�㖄A@U��&�@���]L@��ɠiV�'��� ��F�X`f�q0��@�m~���|2a�t�	�Ond�����pvt�X��B�t�DZ����Q	�r6̐����	��-���?wk�OY���������Ĉu�w�u@�r���&h0B���O�x�	�%��\�#\�N^-iʝq%�������!���Cak������9G����.�J�XL�x�ğvktkG�Y<떪�f���^d���18`L��m|:�S�J�1a^w��yy��&rGVlވ#�D�A����$�g��[o�մ���ƍC�^����<�b�<��/1�Ck3S.��q�h�%O��w��d�aW{�͌��	I���6���������_�{)�m97�^^%D}�+�j�U��/���c�=f�!��W�ċ�������R�$�aZ��I	hI iE�	����+�1;�x%�q��M�L���#A>�����v���3�l�s[�y�H��Hk��#�8����7_7&LV��߿Gș�U��w��F
B	��9m�4�9�q?��Qf޸^*�̸=?/��/��$`70}�~�{�i�1���v�i��[	�l]����>i�)�ɰ��Z����uG�g���(�9��Z]�]׷,�^�����ծ���8��LΤ5L��+��{�a�7-d:��������ә���/j�T�A�O�ϑ�1�B �02kFy1e�5��q-D���	�׽!j������ϟs{u{�1a֎�]��~�j����!Ӟ5�w,�0���
j�@J���\m$�=�`�.F���Xڎ��aFI��/A��#$�|P4T�G�+��Z2�=�uK��O������d3���b۩W�2;���_�u��d�����XU#  ����-"K˻>��I ��</�</#�ԉG;��~(�Y��zU�	�0�	Ԏ������<.�%��\"p$yLS�̡R��5�>f��~��b����h$:y���u+fg�>?�T�K�
#a� ��$��;`�m7Ō/>�������f7B�T��2R��<�
��	�a��<yS�y��J���Ȧ�"?�~�̕��#��PcE��j�	���;`e�x���.�l9��٥^�Ć	��Bgw[�-Hf;�կ�#�*G@ �*������Yl�Iv�'d�
����U��N�{�)��}衇h�5~v�t\�W>(���+�e��~��_��&��A\2"���0U�̚�wx<5%�����ǟڭ �s��̺���UB1(��1d�:�k�=PSW������wA`���0��@%�̙!&|��ݎ@;v�X{���u��-z��yY;����2�H�2 ��բ��Z�.�
��9C��|��~�����׊��� ������,���_u~����X�3���yN����ԕ5�c+ոJY��{t�}��Cɒk��	����,"�u^�{&`�ES��ڣ�I����}���x#���)�-w9���\�`�*�^������U�x,�(�B��[�w�}�8o�O��n��!�F�q x�����(Cpp1AmE�9��E��jIȾ��:Қy��c����K.����_<_��@��&P��(˲��(r�J����VԤ�(�ӈ���C	���x4�I��A��kH�CD�Id���X�C�E#�J:3&�/Z�q%��Ǘ�Rc���{��eW^����9D��k���/���l�%���&&?�0C5S��<�N^�B�����ɱ�qP'��b9u�<����9�8Q-:9p�hx,��j���gxG��+IH�m�13gy�^����]�@�/E�_�-eUE"-���|1`ݏ����4oI~�,�"Q�X{�n�߅ߣ��`��c^����sI����4?Ck����� ����Ngc��M�_� N)��=�e	0���%��!G�|S�6�(,Z����<_�a4�<aw;f���|fT�����r�G.�E�=��C1f���drvQ�UGXT "vJ�7Á�.� k�&����R����m�8��=�<���ѣ�L�����"�'k�æ�,(;�J�!�L �s΋du�]{-$�r�6��@��A�G��C,��T, f�='i�a�)`$�L�5(�R#	�"q���b��/���D��q:�GhN;&�tj�9?R�c(p)?���
,����n1��k% ��Zl��$�Ȝ��;H��.�w8�A_תI,�����ܼ_��.��k��<�ǿk����Y�k3X����k�����>��L�x�zx\���������� �����5�s���9�
�d4��|�o���ᤵ�Gh�&'`�>�(mꚣ���_�y:�&L�`>'1k��X��n˪#(��h��}2
�X���#��$�3=�_�Q�xn���11L��1�U�Ԅ�Q�gFK�H�!��fQ��QU�¨�Fc�-���4�$-B�!x��#L &�gf�2�v7�؊���:������.�IC�&�r����	;.�'�MdO����ۻ���^�߷J�,b����kò    IDATA1ӌ�TD,( d+ˠ+ҝ�n4@�!ϱ���g�%̚=O=���'J�gsK'y��X�A���;ݓ��d>;Hs��4bv>��ܠ��yl?Xݟ�Z�:������E�+pҵ�!�ϼ䑖�������siQ�㦅�MC��B �3>ȋ��z�U��[<��z)�Ō���i�����|K���;����9 ������_�;Z�*1@B��?��dA�ei�iMi���~�ZW=?րa8�ψ��+c��\</}G��~�9�YqQo�~�$LY���y�_���)�L���\�VF]�4ymd��+�?��12��f mR�#�s	�t+6�܂�'�ȧG!Z�DJQD����@8Dd�Æmj^Fޤ���<��� ��:�-(�s�%V8�v]NID&e���������gQO��gpZ�2y,d�l/�#UUg�m���5����>j�QD�,b�,g}�|�bD�A�|�-GȀɎ��A1���$�u��{к�*J1̞3�b�h��	�st��\�߹�k���$WcC�6mP81C�r��g��r��4�Z�3��bx��Km��p�	$C��\2�x�ƼV�u���d���g��|����Q�h:�3c]��bi���,&6-0��ߠ���%	F�6�y]<�����1jc�t��_�9I����6$_,_l�1�$22�Y�׿�u�s����Z/��R3�5F���/�[QQ�L�o�]�$���J\�u1����\���c�g���f˵ 4��q�2(1�:9	²��L9&�I��aj�G���ɖA�-�)Gt?�_���5����H��cH����e��0o�L��7����M0	�d�d�
�֮�3�b�.ԎD;���Ŕ�(��w��9��N��"�Cј�-���nM*���$�!baI�?A�u!�p�B>�agA���l4�d}��]��a�D�%��ېˤQW宭-�-gй<<�G���z������)U\��@W�T~���h�*�G�\�W�'�z�o ǌ��.m¾i��A�����'  �3bt�~��Ѧ�"ޛ������R���6+͛J�Gs��)�S�S����޵�h��f�w	��}�XkbYSX?#�Q&�/���;ǘ����܌8b̫��y�U�r�9
@}k��'�+
��:#���ճ��7�a��w�'��K����l��*�Z��z�x�}�!�����ƨʣ�<���K��DC��嚟�&�{Ձ��ųn�J7���g=�"3�J(9�9k�IMX )-�T^��L�@@9�r����Ap�5(��q��C���~�>''���ٺ�I�'"�DY�ǙjټC2ՓN8���,�����y�GrHF��GX�����&E�"U���G��C�A� ���g�m�H.��]{%��i)p�8�b��G1+���.����)9F�?�	j��y�1�D@����5���O�_ % �=��@Z�����{�b��"y�b�bx�C� 4|KJ��a���MJL�x�t�bX:���Jc�U:�ym�E)psSVKG(�')H�բ׳�����32�}��e��� L f��ƘL�a��/��Ȣb� �0?�Dd�g��dº����>����R!�3�j���H����Ot����";ڀ�1K=W�O@��#1�H$r�����n�#�ַq��5��ѥHj�t��sH��h-��J(�d:�db)(wPj��G@�7?5Ȋ��3M��	[��	�<f< _�^:��qmU
'��X���!(��D��>F���R�H�@8w����W�"����*����ǀ����&j0{N����6c�,���uf�UN����1����K���D��4`91�zeJ�C�����O�e-Mx��򀋭qb��3�$h�Y�(�c�͚�D��1�{qI���6�JYC�$�3�g�'SK����(V� �����3�ߡ�Y�RR�\��`l��DF�y/=R�K�b��d����\��~�z˓���x�rF�=锲$%}h}�F7?K}���63�a(�֒,��7�	��#AX�Cf}#2e�u@X���!ه��¼VE�p�@+�����z��X5�-��{�UVI�M��'vo�9�	�
s�)=���9�	�YR[��<a������;b�S�����0�]�L����vP���|M�Mz��vYǜ]�xf���֣�͵����5�Oŀ|R���E�0�m��wA��;s:��F�(
�8r�v �}dP$k���9���;��ڌ�:gfs4��"�ܽ���J(Q�F�C�z��ۏ�������q�@I��u�x�g3>�3}K7�Gm
��٬ed��0rYT���1����v0�e1b�9��tJ���'k����u7���6b���X4[� ���,�5p1hް+�*IKڈb�� t����dN�\�!��y)j@�7��	�f.V�{�Kf�Sg	�Z�҅+Mf�:5S��� ���6TW��*�z��n$6��9�Pda�Mv&���̈� O<��������W����xɊd�e"�2���j`�0&k��W]uUG%2����,��{d��X����ؖ,bޓ�
��0a~VdClT2�oai�hu�)ʗ/���z�Y�֗|�o>i�����]���~���lp�E3o�˷�	3�@XrS����v�x����Â�l3q�0���C]*@�Ў�X4�S�ZQQhkrR�̲� -�56����꾨oX�d҅ �-�-�݄L��h2���3�dA,�W۸HG_A���=)sđ�߷�*W_m)�A����j������'�����Ҏ���(����!�T}�r�T���͆�[v��MNV�z!� N�H��1c�
{~I�P1�
�z�.�b���A'3W��En<b6��8�`Դ�V���E2�� ɾ�D-�gs��|-�s��&��Z�~��YM�m,0Es��O�\9En�ǝD�����;��$�Bi���"�K a>�L��=��ö��6�(#q��Ŧ۳�Ɯ��ᕱ�}�	���4$x�R>[�6
E#�|�w�H�R�u=̲*�3j4��a��>�|�$��lvQ���0:�@�M�ϔ��b�e͊l�֌��"l�IW��V��/�7�,DD�'��}���ϜT�k�b¥0�D�A�(��A��e3EuU-�%uУ�?���H�J��H�rX4�sZQ�(��m�D�\!�=��C�G��ꋆ�� ��H�c��p!n��f��-b�bQ���؋ǋa��ߣ5)d�Z�7Q�z8����t�*M�|�Y1`�Ǥ>�|n}�,nnǀ�^hY��h�X�HU��WU,�����"[4�|��OF��� �����R\�t��i��1�`�c~�,�)�2�|�B�&�P�! H_��%'��㎎��iI ���L�U�L��uP�%8��әK��7�LXlI�?+�t��zv\�L���f]Ǟ�B��g��ڷ�$���<�A	u����l��{��A���� ��mDt�K�|#� S~��6��$KE�	�L��%]��Ra������ޞAX�`�6�bǝw����0;X�`��'�F*)�Q�����t�k���. WFW�� ���u����n-eI&�k����r���'�0�Z�ԆY������^=q�1G����@8^hÒ��5�G2Z@�o��٣c/��(��#F��xOdKI|1n�<	-�f$���������K�!�Q �Hզ��V�������=� �4�d�z��"U��d�C��G>����q�K/�1S@CMo,X� A,�h2@��|ɠ��ȡ�6)Wys����Y��-�J"��$)�D$h�*١X�LaE H�g�"��Tr��tlNx�:�E�����@�lS�"8x���#��1|���^���f>ٰ6 9}V �}�Ii�78I�E	Ѻa�[o�m�#uM%�܎��JX�F��f�=0hض(ī�s��{��A�A8D*��Ի��{o���C�TD!�6&�.R����PʛdUcq	�	l�Ŗ5f4���s����'v��|�F1V�JS��,	��P�Ed,O^&\	�����lwY��}"�췒i/���~��ğ��8wR�c���4&L.�6�:���%�ƀ~8��г�B�b+Z�A�e!⥬1������0̣�h,�S
jM�F�~��C.Z�s�b򔻱�y1��q��gMPR`̲ix�� D)(!oi��tc��>m9$��PM�:,!��S���P�GQ����x�g硵��d=7��\�R�����L{�@cƬO0�� �"$�e�E�i�I��h��?���xb�2��td�<.����c�]���`0=�%���RkQ��x겼F��S��xV�"�&`�$XW:_�=�`��tA����w�I7"t�^�9bz��kT%Sv��=�gϺ�&YK��JƐ�ŰU����2��8���=_���{�m�Y�m?3���G�rS�q�ؒ-۸C�B	�I @�!���mll�d�@(!(�dzI���EN�Ќn�V���g�������[�7�JG���^K:��=3{�-�{?�S�(�jT���$Km0j��;�i���[�����)�T�6��[��p�H��Y�Ѧ�����g�b]r���P4^i��h)��D��d��[�uB�u���2�� ��2��Xnx�b@��k�yӲFG������i�*�:�vڭ�W��s֟e�}=[�	��Qk�LYbL��U�ȲV�*�)���s��Q�������f^�<�ݣcv۷o�Fc�z��g��LN9[ъ�J#�f�Yg���bv�،��Wm�=�b�i���k[�8�Vֲ�8��Z���������3h�S-�F����6�w����A��G[Pl	�n#�G@��U�d�3'�z@C��rm9�4��A?�Ctar#t����hRć�#�ع&Z,q�8��Jb`�S ��B�)E:�9F;8������(L�}Ӗ�V��`'���g�� ?0�,0a��jZ��n3I���m�IgYr��7�1��-+l��JT5k�����'-{�v���oي<�z�9�U䈢�*�~@�RK: \���䣟d���lk6ˆ�d'���|���W�򕞶���G:0񼴷�a�ݖY7��!_Ch�u����1Wh���/��l��B�|0WB���8�p�Y��n��5�-�Yy�~kc�Y�6�Y���L��t�1*'�3Nw]V,��-'\Ӱ�����3]��ZM�R��d �d�֎�Z1!�����۱3��܊�=�vD�� Hcڦ�Bt�U��HR��+�?{�:�o����,�;8;�-b{ۭ���N���;�� D��Г,Sق(�Pk`
���h���*�H:3��}J(@b ��������
`ܔ+�a���(��)����a�Jq3���M�B�V�ݚ0���=�^��ㅯ!�o�z!=7��g���C�����$ɭ�6����R�X}��x��O:�F+��N��.�D@Q�(m[�N�l¢��nw~�VYfլe��3a䈘�R���zo�j��ѶV#��Zݝ�ĭ���XgUl�pᢧ�(����i;���B�*ڡpt�cN�7[�/6��~.�\���^���΄	Q[�}��_d���*hmIl��?�f�Ǌ��Da�y�H�(v�H�R-�E�7��DY�'����L�u3��jQ�|��#�05<|$|�����XEX��]vb��Y�=y來��l7��6�YEC�]S�Z���^9l��%vOOb�굶s|����h6�T��λ��{���#�p<@IX ��*��2ay�(̯�7��	��pi�������*��sТU�[�\�ܫ��Z(X8�)�DV2!ll�%�P����c�=�x�M�h+ŢsM�?2Lx� $wռ����m�1e�(�f޲��^Kk6�w����*ǜbc�A�`���|D����ylڶ�ل%?�7���;�*ʭ�6�ؔ�@��U�"�u��Z�8��k7���h�V�pPJ꡽�H>�l�E�Z�X��������ąLx6P�n���ƈ�,#c�s��m�4�r&�_��w&��*M�1�8H �JR-k����{�e��A���L���DE��Jkd�W ���L�[9[掙��s^l$
S�xm�E=l��;)��I#��rb��Yê��f&XےV��%�Ț�������M�׬���S^��E�Iu0�T���������1v����Ģ>�X&�H)��b�ۉj"t�AP;���0����~Z�q �$�0^U��>�~Ђq��P�ó�F�@E�1E^���LZ (|�@ AX��3�p��IN`�y�驤XSN�p(�~�?�Y~���
�iN�L�p�n���F���;��;�b@8�f�j�[W�9�@)��M;,����̏�k+Y��/�ʢ(6v�a�FMw�E�;D K��$�Z��l,����Z	�G8�e���(Е�p  <���3�X�@k܆��{A*A���|�;ߴ~���K����}��lot�����=zzk�6C�Ll��aI5�v���bbk2���H0A�x�Ҥ�t:�I���8K����7e 1��/ ��F��bma,�B�Q�g����N�%xiB�Q������#�2��ʽ����,.7 �m�V���p��y .�//�<�xFb�7���qd�8��$���#v�Lj�b����641i�ֲUa�7�'�nq���m]�Ҿ>��ݽUk�$����ε������w�i���@'��{r	��")�[��_K�l�?l��
�(YCq���tb")���&�⌹&�Z��(B_J�XA�@k��8�c��rM ��"3���9' V�c�.����yV:9��]�Ŝ��z��"���r��s: <>1j	�0��hV�]�j;��-;���[#!�0r���"����#�~�&���3ូe��I�Va������=:ك�� B�<=ȭ���hi�b�J��M�҂$�J'�g���CR\C����!g>�J��`J�	�G����u�	VI�48�8�q�g����3g$_��$�ʢ(���W_��e��󪧮ڽsc}rt�(;k��d�U��i���� �9kPiL�T��=��T:���PcQ��������I�p���|抛�(�,Ei�����\��+C�<.0-�u0�D^����ck�2S	05�`_��L,C;�K������+>i�+^]�ZϮ���ɦ������)[1=i})Y�5K���"P뵑�j[�ٿ��vgod��56�hYk
�m���A��������1��O��b�J &}�s���9C_P�A@XrD��uX'ז<!ǜ��ø���}#9���o��J�a�B
��@Mǜ����M9���&�x��yf��*�IG�� |��g��������y��Ƭ�vTV�aϾ��Gg�!�b�UXЋ�9���r��|��;�a�w�����YA�R��m�3_�԰�,C+d��� S��?~�l�+Q�#�t�<�,|���|�����2q 2.�����bb���"s�EZ a�2<��5TIN�͵��+�w��qM�cT�L� PO�37�|�O>��=Ky�y������ؽe㊬qN��0vֈ��5��&�њ���!;�<`g�X7!���r?���`N��w�k���^��luM]O�Nb;4��ϺW�����S������ߙ�Ej(N�"5����e��bLg��'~��LlX	&3�h�L-A���Ľ�!Qɬe6\1��kϜl؉��Sǧluc��r���qݲ4�
��R����=X��=�5KW���f��F�z*U��11:fqT�;����n�>icͻ԰e�#0py���{��/�jCK��`<�s��ń2�=d�jG}�~���u
�	b� �r�s�	k�Q<2 ��&��Zs�ZLx)Z�Ϊ眹��䞞>K�G4��k��7�m�ն��Z�l�>h≉� B�*x[Lzs�ik�qK������_�a�+B    IDAT:ά�Lx���.�
��y�c�ѕ�(�q���\"�]�2���L�tiG�!]Gc8�e����g��RҖ�<�'��3���G��0Bf#�r��ƪ+�xU�6,��kHW"��-�c� ��`�9�.Ϫ�'�_Z��o-+��Ʒ<}�ևoYg�4[3��*mt��ƛ�6�r�w�8��}��	D�p��aC�J(�W�dV0������En>��shl�I��ƕ'�c�NM8�����:&�âZ���2��yf5�s-�w�Ee�����8�/@�-k��������<�j�bY��n6�Iw@�՛X�J��C1j�6�vB���	[9M_��Yw�fy�I�j���j�eՐ}�?���m�g��pD��(���^�!;K#��]w�=�����!��Ć���;��X`X�'lsZ:�"#�%-�0�r����s/��:�/9��o�y��&�D�$��!˓#�+:Bm��<����WY:�p�U+�r�M�ŝ��l��$���yVԥ��=QݶWW��g�o���6�5��}�0�p��r&����6v׷mMlVO�	�V�p��I�ZRK<��,I��9B�/fZ��j8�$H,�I����T���F�2��!��31z��1NȘ�KV�|f,���
��(8¸;t,Ϣ�x��1a�; ��8�.�A���1w�7��ۧ�z��B�~>/�Wmߺq�=s6�%Ӫ)�vf���ο�v��s<�3�"N:_� �י�Hc0�y��MHb8:^�N ��_�r_� 0�I�ɤB��%��ΗY�Ux�FaPc��i� �@z��ib|��ꕒ�Y��u ` 0�zp��9���{ՙ�0/t0IRL!�D=P���P�E�q�Z�e���(�ά��6����q��N�b;zt�V����ܹ7��"u��V�j#q����G��p����nzl)1�+�\~ ����羻|��.3�A�5�e�p�$=�A�R&�,�V�VR���h�0i~�@!�HÄ�@Ӷ���9�c! sK�~�P�8TB	Yk��X�@DdA�SCLXKOq�L`b��)��n�f�Ln����B�Z�z�e͆ō�����ڨUmGm��~�y�>�D��;�x����<ށZH������6qwᘫ�g<:u)��@f#���d��#3>oD���n���]�նZ��8u��\%iHㆶ
��5O��c��}�o_��/~���\���}�+_��~����N�*���T����¤.R�T$���*�B�,�|��jn�xd���7�p��.+?��o�ڑG6V���'���i�0L��S��_~�m|t���>/����>���19�ƈ��Y��>`U�+�6(c/zы�)��G��e�]�E]�������*3J%�h4�<��I^�:#�2׿�,*?�9l�� ���֜�4K�V�&�jN�X��
Ḻϕ܁עj'�|�#�^�Ɏ�[���n�z�)�@A�Z�;J(��<@��8��Jl��{�Ln��96i�hR|���fI'�8��Zݶ��m�����F��A�k�SO_�;����B���N�Lfm��b���e *���{���߀%�(*|M�H *G�E�����9��9��7,,-Қ�_�V&�駟�u�x|�,&l��(�M ��ϸw@�	��Z���!'�8�:���d��C�Y�6rWR$k G��i�*��k5��-����xT��a[s�k��X��P��RƓWHB��2[�OYv���]�)@8���̤3�F;wn7��q*�t�Z�f��Z�W�#���!�VO[sjW����_���ojk��f����ox�k� -5G Vj���L����m޼�ﻛ ҟl��6i�3@��f�ݒ��?�	x^���Y�X�p�e��n��e�5����[��
��v�QG���?r���w��o-��{;,��W?5�UޏI�C���(���(]��X�^���yN;�E4>�b&�����B���U0�7�Zq�p�6B�2�bxp��^�[�j��֌բ�Fwo�tf�z��5S�	(N��׏�#��_�j�U{V�>s�nY\�ѱ	V�zO�)�ӍbK���8d�,��
�+�<ڵ۞2cvR�׎�lZ}|�b�����H4-gq���ց��f2������Bz{|_;j�o������% ���X��i����l8F82���Ԏ��+��\e�J_�0�BU��b.���{ca��6kr��z�#��Jh�,�b9>a���l �ǜ�qó;#$��i�B�pʚyX�ӟq��F�аM�O�Ӭ(�Z�I�؞dȎ:�\��z�M��m
*��E�G�,JS�6m�w�n{��^'� \DG����r멱04,�&V���i��}���<��x6��H��L��]N�l�7~�7|�-��E�J@ZEj�[,��_z�.�^1�A�w�ĩ�'`c��������Y0CkJV��Kƍ�+�2�@̳R���"�Jy�EѦ���=oYv^���[VX�l�S��s�s�=�%��w��_���Y���		�0��L+���xp@g
��AC2�1���a�����}��C��9��h����Š��`>��a�l�]z��G���/�'���&���q�͌�X_5���������C�En��cK�VZ�w��9�ҨϲJ�mٺ��vl��`ș�4�d� �}a@ވ�	��;fϬ���k���������ӹ��"���Jl�(��������^m;v�q�kR;��f�w//L�'֣	"�U�}'���[d�hb��É&&$`���'��	�д-�v�0�K��5fd��J�P�eq]�h!���a|1>���&���Ҹ!I�()|d^����p�96^�hj�8��{��W�cםg���)���L�2�"�-�2�[v�7��v��CF�JɄ��[����'���S�̼��I��r���g{�lUʣ�� J �:�SI��A������O(,���bA�ve�/��kQ`�,���2!�n�G�w��#����y�+�����uñ/i�-��<��[n�ſ;��Zqo��޺� �&�r�#W歳(̀���+m`u�}�;���W��a��d����Lh|4���Я�6��)��P��.�*�'�U��?�4���ц��|zp̙��:�T�V%޹�Y++6���^i�}��OY_���b���ZV#<��"��`E�,i�YT�V�g���6t�S�	�}�m�۴i�kp}�U?�A�>��ĥ�I8{ r#ʭ��cy�i�Ql�񫯲��,I3�խ�h�C��FaS��Ib?ٺ�>�7_�Q�SkuOÆ�T������r�䢋��O����ov�e�+>@S&?�$&JOz˖�v�Z5!�N�<���Pp=��U_jr�R�0��~ ���|.0��%	�����31D{hR
�%o�����H��zv�AD�_��0{�|��S�*���l�ն.��N9�,�)� �@�"k٪,��އ�����o��ﱆR�0�"�O��S�b�؉	vN<�?��Y������7�f.���~�ɳ�|��ޞ�J�ô/ɋ7ݏ@=��5��7J�^y�΀a���W� _|����Ӯ3|���4��}��?A�+-6�2��"b9���X�`��?g�@�Y�J*�[n|���� L��ac[7�&F�A�t�;�^��+m��#��;~�����(:����3(L7U�X��ѐ8�ІE�FD�{��^��0� ����]t�ׇ����+71�@b&ZqC����o�Z'�b���H���׾�56�_��9a�q�vo�w[o԰zJ�Vj-*�Q!")UL�v\���[uh��}�5}��^{x�N���M���E,1��AQ��zl�G��qbc���]��W�ꕫ��V�p_m�\�E�-����s���s_��MLO���a��ٕ!q�6��"��9���?�R�ir1�Y@5�Hb�$��N���`�i	`��@��� �P؟�����LL@���/�R��f�x���*$�iBr�7�����P�ǽh�`�`�!��E@4S�5�,��Tg�����}bi��.���l��ô�
Ql��X�S�ǿ������bl�n���.��-X|faYF\w!�M8&^�s�C��������r) �͸a�9�?2�{ �ō>`<�7�^��=��p���M>%�@�s�0�9xE8.��x�,li!4�j喛��ۖ�׌nEv&c�Y�<�^���m߻�v�O��-�='��	;
C�ԑ|���ʢ�����'?�4�������C����װ㗼�%�z�������WZ�
�I� �k_w���,jOZ_Դ�[���3�,oY���WN����.�78�i֎�����m㭛mz.kΖ �a�Ԟ-ct�I�{ѡQ��e/��׮-*��5o�^ �ÌjUkf�=�Ӈ���w�w|�������0��OHL@&b�F���߀_ ,p-ڭH�`p�4%��Ľ�ó^��	�Ra.��0����ώ]+�HzF]G��k3I s�0�j�r4�Pa�R�`�O���-a#���cR}�A�>i�ܷ&9@����������j��6�(,��Ͽ��F��`X����	5qa*;[����}�KvםŶS|�K!!x��$��\ �yC�Qʲ[�AX}�O1ae>���L�s���H�ā�ik�,������Ɲ�7c#S�`���i�a<�	��5|�w3oX�q�M�ZZ�$���׽{y�0s�[޴*J�z�}v�ΰ�/��~t������Z��0/V,4��ix
@�B+6�0 h:�������h<4�0e�yp&:�R�Ť�o
KÀ<ڠ�-��R��e��j'�NF;0�g���W��@ݬ1a}����齖M���j��r�mO)�=��Mm�aFT��/v[>�ֈ������#�3�.G(O$�lM����	�31�/8�<[�r�O�Z\+��)Mo�x5Ҷm۹�n���695U��E������	�~'�|��4O7(3��7���a��'&$읶���/Vǳq-�$\[{d�v����=�هLD�Tߊ� ��������sM�	��XV���Ua���!2�CV��@ L��D���}�z�^CB �~�m�u*���*#�������I�:ŭ
^$���ʨ�<���۾ioy���2�C�`6f�O1aL�n�%��d.�{@��B9��º�����M>!��,�ZHO�Ї܊�8=;�#9��4Db��z����g�a�ϸg�k����/
�ݺ}���fd��w����6,_��#�<�ЦU�n�iLu@��+.�0��V`1at~W�Q8x�O|��	 k�Ya	�E`R���/v�ba1���\@��]8K�9�8����u���V�,jLXo���	WҦ�F�+��<59��F��_���Ҹ�ޱ�6}�3%Sͪ��@��͂	�l���SE�U+�}�+
Lګ�� �9,j�T
5���ωC�V�l=�pk��*q��Ԏ\SN�d����3�8Ma�:`T&c��,_z):.\��59��2F�L��Ư��1�c���Ɛ@T��1S����!��$�;iC�_1M}�x�Ox_YWb��a|b��O	-D��g��j��	Ÿ2&t�.��-��νV��-C�_	w[V�H���ń�����aڌ���:Y�a�� �d\ >K�v�%k��
4��|�!t|���j/@�fQ�V|/�@���c�nYv>��p�ѣ�l���l ��pʱ'��_�2�#��.�?ǔ�I��!�#@�ae�sF�&���ԧ>�lW&.ǱZ��ot�x��������W���>A?򑏸�,P�х �s9�y��)X�<4�o�{�ڪ�ׄ{��3a4as��Äٷ���គ�c.��n����mőO��#;v��[?�ż)��p�	�Lt��� �Yy�Y�t~�@���s\j�r^4�g\s�]p�|�l9�rϚ�j��ݤ���`j�#�qM�E}*kF�mh���� �q�Z�E
�C���|��o�/���5���u���$����p����I�P��2?�ǋ���g�M]HZ�
��X�0�Xp��pұ�R"U��+3]V���@x�L�@@X}���0a����|��@D% �<#�'�g8�y�(EhgA�|<�5\�4� 9c69B�E�!�q��!�@(G�yފ���_w�ۗU����wl����+��1k�d�yͫ��[�{?�ow̱Zs�au�&��V"����F 5zaj����@f%�-˩�b���qڠ��Z�tP>+�+��a��q���Wmh��)뭴lǖ�,)@��o�ʆ�"��� 4r� �n=��Ӭ���D�u��u�glz� 5��o8��{ͤSYɒ��{�ܑ操h�>~�E���K'���U��W�(4dXb���sorӳ0����Ҁ;�rɆ�������^}�1��NOw�:�Ȕ���p�$	z-�2C��!h3f����P:�:z6@͙f�8$���P���"8� ѢP��]G���i�Lu"��!)��j�7�T���(U4bҘ���q�X��E;������4a->r��Mń���&y?�#�����4a-���M=����N�ue�9�܀#֢ȹC�~%>WʱH
 ��S�� i���p� �D��=�E�d�j�z˲���+޲y���%D��=C��W��z�k�����5�a�@�ۈF��Qd:��P��TMڏwS��u�Nۮ5��q<l�kʘ�M@ŵ�4[r��pֲ��~{��^cCu���V�R�������Z-J���A#1�%�=�Ȟ�,�)�^���a�ꈧZ�j�Zݶ���L� �g�h�ζJ��:@�v"�j[S��平&K�X�5Q	.c��}�q1MڃDwv� �C"C;�m!���dR��@N]�),g��_��~
� B�T��7�K'��hu�"#6%G��s����X��� 8�F�PH�>K��؇7��ߴ�X��D@���;�̘�Á^�<"����zO����e5�m	������3��� X�c.4�Ŧ�A����|�#ǜ@X�,
]{� ��[__gh�n�ǰ/%)��V������lN.�u����P��~�2qÅ����>��4M�7�x�[���O���C�����t 4�f�yϻ�.�������'k���e�,/nN�U7@� 4���̀&��<MT~�L���|Ql�L��W���Nȑ:[����V���?蓂���<�.��|{�S��;ئ�I�ڻ�c7L�R�<|�)\���Fq͒Z�E�~[uؓ��/{��s��w�u��~�h��v�ffx�a@T��$|��#T�M �-)����ZB�u2���\���y�P:'dܳ�е:��s��_��^/��K�!����Z����Y��X�B��sHz��bބ㑬:K�`�ra^J:�3@�^�x�����U�_h�.�M
g�B$��H�S"��o@����c �*�\��9�ƊC�6`�UeG�\IE�0E���A��_�Ӑߡ,�馛n�j�Ax�O7�Ό#GD��TQ;��g�%�t��{����;;���sS�):A+4��F6��j�@k�db<�[���T��*���H����>����B ��Ť݉�ʊ]*�w<I����nN[N	 1kY�R8S�{.�+�����Ψ��Z;K�V�əF�h�P����1E=� �uO�0���J�G.y���o���ŒP�����<��7N��~ ��|-|�\�o#��ZES.����4�	���_$:��%�%q��x���g�TVQ!��3��z��\t�ԅ�d_�H��/D551}q�N��L1S�E�EDa��3�2)e=��+W�k�cX�<#�O.T֕�E�7�����e-�^�w�����s��{�����U����֝b�^~�mߺ����d�bt;*$�����y���`�$|�< �)�H���f(z��>�1�
�g�h5J�����&���)_���l�AW~�`    IDAT�d����j������JU����b��)Oi��B�����1�Ez�I͊�d�N4ݟ����췀S����r~��&�;�ׇ��������Z~��@�쁞?_�?>+,����H����^���C e�IǗ�S@�q�����G��F-0���_j�b��f�V� �A��3��y�	��_��_v���)A�$~!�D��z�~$e*� قci^�K8���H!�'B��k���S�_�� ·�����ea��_�{��3��R� M8����	§�r����}���ǃ�)�W�It,l��A��8�b`��e����ωF���O�,2������ � (�=��P9w:�
��^Zi��%[8QO�}�<5�C�e�d�:�_�}���iR g� �׃vH�E����g��dL����u�`;b:� �{|vG�(�н�K a�L����?t��h���<�s���s��/����|����)��s5�B��W��.�[> �:�^�+�� E�=
�7rȨ%;Y��U|HDE��983'e�s����j����M%9���sN�#����i'ji!LӂT�1w�5�\�;g�yfQ�j��y�	;��~�P{fC�5ת=.GP_��5�~�Q���s�SN�`����U$��A��4
� N
'��F�q��ly�a�46���פ���~�������=��"��wz��4
����=e�I��*kC{s�����Yg��"[V[����)}0��m�`�Ԙ��n�b����� \<�����QW �>&�;&٣��r�	;_݈E��C��X�a怀Q��T�m�C�C�P�_�'s��v�ii�w��4����&���,���Y0V�b?���|���T� �H�BG� ϊ�8cpGa�r�GH�X�+"4��p���:�)�~P@x�����ҙeI���@��Ɔeնo8<��AX���(L�7�,K����1JĔ�C�`�rX����Z�ل�:�94���C������i�-d��oy�T�V��L3��)w�%X+��v �b�{^x�=�+���
zSP��3 �`,>��q�k=tt2i��7T��ھ. `>J��ޢ�K()�ό������<O����y���@X��,kS�$cO&{�a���V�I|̓Ї�9�<�$�9;[�-L����-���:\,n�Lt^x�����l->
���/JI��K ��C)�R���s�vl���t�<��O��]���eg����4М:�ZK��L����#���# �f��:�02�r��� ��G���W�)�Rv��,�.	 �zj�)�� �`�P�J@)�X��\��xY��öju׆�S�ʫP�����͢�O���J�I��;�*k(��������-��d('�&��i'C�ܩYϠ�JY:KgW�y����`0����"x0�m�k��[���~�Y�k��֣#gB�f��s�CPS"�%�N���;�$tg�q�:��clUa���w�+ic!'�AH��W_�q *�P�x�F����|� ý��k.�� ��Y`�V(�
CS vpK�=�Vj��<��������:�n�kL<7���w�(k6����^kΰ�4���*�m�i:��������H���@�@N=u�_ܯ)yL9&�]ך��\۵ȣ<`-�+O�(Aد�2��������F��)���:c`�e/!YDphq�-h\�-�/�z6քS�5��ɚ���kM�\k�I�x�n��~ޅ@b��Y~���х�ʅw��ShZ7!q?F�-T/�c���V��\Q��0T�g%��:�LXm�X�:�[ S�B1�Pn��h�\.�2,�S�V�d����"<�,�k��J��x��#��d"��)�
���kkY�������5;�nn�<9B�y1�=��|p_��lN@��Z!�٭�vj�e� u\��l:�R��_;OMݹ�N�n�u�ɱ�{�u��E�t���@��������r����5�">��н`jᙏHB	�ٚ�\��	�J9����hC��)� Kh����Gֵ�g;t�8��n�� ԭ�@�����T�� ̖��\s͛��	�����z�C���3�/Ą���k�-t�RL�C�Pj�'V�5�Ckx.��^;�����>Gy�X&\�T>{��W�� ����ڍ��U�L:��"���֥�n�^��r�C�j�C-��jEO��s���BdO�5�nv<_��:I��]{�o:�3v.����?����U��mj�\81���\�B��9���>t̡8�O�Av!@},�.�J��k���7� \*���U$���5��n��bq!yb1�8t̡8�O��Ɠ�������#� ����Aᕻ��2�:����l���2�����x\��C�j�C-���c)g.Ĥg#��ß;�r�� <��vk-!�.���5�!Mx)C�б�Z������n�Z�.�Z�Ơŀ}x�0C7I��_{�o\V9�舵;��35vA�'TMLZԂ�X3���D���d��nN�<�VP��UP�c�����	���-�U%I�|�z��}��Đ'�P\���L�ӱ9�%jf���ۻ�W�����Sx�f��y�����w�p�({��4�J;����u]�s���m�v;���<݁F/i�+����Z܇>���ؗ�Z$�����X��<%�h�������V8ǦiJ��篹�7.ktsk~pc�����6����ay�0����w	h�:;'(B�1��<��=kH���X�Ұd�i�p���� �G��8O�ε�����jd�a������S�49B���Q���I��2E��$J�����!lS��HR�}j�nֱ��:�¸P�(G�����*�	STM���+m��?�P�z�i���3�ɭ�.k��'�ND��Ͼ��|Ӳ��\�cۦ��q�AiF���3���yl5�ޥ�Q���\@W�Ȁ$����	�_����Tǆ)�4�R�<�&F����C��Ɂ0���r63.�䳁����ͬT} �0�N-c���Rjm7�	t�b��\��Z���|L����3��c�2�4�*L�Vv,��wҭ��®�WY�*��(�X5�9�td!/��|�6����иA(�!���~�0{�� <q�EY�VD���KYR����P��njS.��ԏ��7LcQ���q_�ܥ���k�K��򷵚u�
���TUb����m.���}���w��!����R��{������)�R�J8�BY��e�،,�pﱥ����X��݄�6`Nt��`57���X�Z���2a6V��v<P&���*�V���9,F��z/Q�)T$i�e�$�Q;�RQ0��ƠԢ ����UyOڳ�:[�eY�$��馛޼������9f���[�ugsa/e	�5��&\Mjv�	'y�3�+�h�Q���:p�S)e,yHm����:�i�IA �F����W\��Qb�F���O�a�}�3X~Q�	'�lZ�B�;�.!�����􋙨2�Y�a23�AX ���,Qas��i=�PLU����'��)|ń�
�<,��f-��+sB�E0lc��B�R��\����s�����t[=(�h\h�ƾ�����,p��z�v䡶�dRmH�ߜ/��a�����K.q�e)i�7�|�o-+����{��-mN"��f�3�4m{���/�~�g�����������F�K=8�9پ���x0X�W+KI��^��Wzaw�
�u��h��?��?�5!l^TB�^l��"�ʂ�	�Xf,p R45��-�P��<��� �S�Zf����*D�E�� I�~�U�:;Gk�w��$�¶�%2�(��%�} ��Rd�g�x�>v�ئ��`��!�9q�I��/��S�}˖-N� �b�c�	
�����n�+�qmI����R�禛n��e�ön�4؜��eq��5�v�e�k��ēO����η�Gn�X; ̍�TXj��P����#O�` �V&�����~�zc�e���0c���a0����9�r<�
����O�	=׽w�2Q�Ye�a��	���4������K���^ĀB=����c�'�"+�;�B@���b��H��ؖ���v�0�  aɀn���l�k(��K�K�'�`�<'8"�J�jW9� i��9��]��0hD[i�����Gb� �oj�K,�v	¿�� |�o^���M���Rl�C�ZGv�i��/�ܲvn<��x���29U�Rab�00d�*�.+<��/~�M/��<�����њ�~ɁƋ�n�wgl7�=��-e��e-N�(*�jgb��ahW/�ζ�8���Ga䅊sk[�wo�7��"�p_1���bcQ�����W���Q�Z�F�� ����9�m�v3"iv2��eIKܩX?_�I��g�1t�! L��"�0��7�W��fN!��ga�Ȭ ����Q�I[�I��֡���6\��5{�o���k1��"a�C;�l`�!��De�7��,���� �]t�c��,���.�j�	8H��l��?��[c��ҡ�<o�q|��7�������9/� y>��ڵ��K_�[�z����?��[������&+�#�ѓ���D������V/�3Iit��Fg�O9���/������c����ڹ�^���l7,Kؠ(�8�,ɫS'9N,�k�N�V��_�E��/F��,�V��hP��;)�^l���Y��>�������J�e��[�1ױѴ�Z���zll�iQ��r�FjOY���le688�+8���B�Q&S���;��X� �U̖��3������|��*}�]R�F��u�O9>�n��\�(��Śb5�0��{-{��?V��BKAE�`xX~�0m.F�lS�������}!?	�ɑ��o 5��O�=�k�����~�U<����E�����pa]*s.;���u�s��8������}C����|�+�|����d�&�gc4 T_�9�[q��
sN>�dg����q=��q��c��o�j�A��m��	;W��k��֝e�{��ܽ���~���*6�,�]���[f+���I�1!Y��h�dx(�>�����4 �\���x�w��M��{��^�A 4�Y8:"��͞�YO�~B�z6�h�������f��a��Z�����e6lY�kI\3��i�a�5��a�Yb�%Va�O���l�;.ge�b����Gj'��am�f�eyϰ�6sKz��m��3V�V��L-����me�ϵ�a�X��ڛ�u���y��Ō$7	D���x�ٖ��arL46�\�������w�f��ª�������Ҕ!&��K.�ĉ�fѣ?'�����I���/�r�s.s�c�$,��ER���/Ӿ[c^�G[0v���7� �@���`�� ��	�8�GO�,#k�~9W�5I"�"��M�[`�ӱC�g?�Y�GinEQԊ�x�7���SO=ud����6��8��<�ЦYk{��f`�����?m��v�~Ӧ'g|�L^�'l�':�	��ɁHs�I'������}��a�	X���Vt�� bP�����X��Ă�[y�jQ��<��x��8q�L:I(l�Z֞�a��ڶ�/����G�bGyӲxڢ�U���ȗ��;9�EHiɄ�J�;�K�]�YT+wp�,NSk�UK����F4dI��%�j��Q{�I��'��| �PA�.E�ȡ!�L:$MS�R%�cذa�O\,��ǒ�<�����k��a�/"�"�gԜa�/�C&.��s�)M�A��4a���:�|ļ��gø�a��Q����a�.spbΪ��	�L 9N}"�N?�tw�}���������5�\�D?c�FB��� �Cb�8�5H m#�!��̡{�<�c�����]�& |�5׼���~��e�y�sS�3����f�x��m�5f߸�߭VA̮�ꊼ�nv�VEn�P2�:O��@`�������?��yq ��
�x=�Cg3�B��x���0{�r׮7�*���XiIT)w��,�&�'��<֞s�����tݢ�bI��X\mZ�'���w�d�	}cP�� �Q,X9{����\��l��&����V����rа�9�k�������oج�Y� Xd,�tJ@�6�G�,Ą������A{k��<y�e"��_�җ<tJ`�6 �r�).p�o~��@g�}�?; Ä5��k@�� uM�����jC9 ��cN��\r�ƽ��Z �|G�N��W��Ua2��|��׿��w�
�q��	'�`�_~yg�^���9���'�"�n���e�6����9����	(�T;��L𓍇_��W��iG�{L��5��`�sЀ5Ƙ[�c�e��������V�Z�Ե�^�{�
�a�p�^q>�����Ͽ��z��y��=c��o��v\�E�C�����n'��X��:�,w�}�_p@�e aJ��c�a�p [@����$Q�\�.�b�f��Ȧ�Ik�T���m��
���X%���l������c�lz�NK'
�7A��,�iY�`Ū�Ŷ���<~�[�ю����۶�ڝc҈ݛ娋͢�5�A�6�o���-�eo͒��f�8lV3��C���x~&m*�!dG�i���g�s�1�MXk)�MLv �2�9�Iʀ���w0Pq��9��#�}^���o�������	�L�߹��s~@X���Ó�1��&���#X��� E�m�{X�|�V�d9���-&�pB���SR	�ym�� 2t LX�ĵ�8�3�]v�[ь�?��?��(9N>(�	��/~�k��E�v΃ �lն�Ap��6�m�G`Hj��ԧlb���J��'�s��o_V9^�{Ǧ���s�� c���^l�}�y����۶<�S�Z���+��C�0aq ����!�����eT�kݺu��7���$�$���4 �Xߩ pX��l²Jd�z�=�����ZOo��m�Ѵ�c�p�����Ǝ�Vi�]�h5'-%���e}+�ĖEm�-�=��� ��P�x� a�$��u�2��5sL�Ul:^a3=O����f��Y;^m֬����Ծ�w_qYFN-|b�1a&&�����ĵCY)���B��cp"-�ޘ��������W��c]ˮ�5���������7��#cx� ,тL���1��$'�m��r�s�m�	�9b�!�s>}���w+����˄�L��/���}z��9c��b���+�饗:s_�YI�	$M���h���cq��8H#��c�>>�<o�qr����o۰aÞ�X[���>y��G64��E&*��u���_d���o�O~��U��E�1�r��蚼2_���,ei|��4�-���%F������J�ַ��l���R#�CL�*+W|��
p-�Y�ֶ,�,�*����v�ŗ���g-��m0�a���,�u�ٞ]MU,��Fl�hOZ�3c����-�"l� ��ٝ� a�+�S�*�-ɩ��g�����E=6��ht����Y���hX-��*�c�6����_g���X�&�b�0Z;�-�`��F�H�?�2���!ib��hh�qMm)�?�'V�&�R���X��Zlh'_����Br����Tp b.(K�$�D�Lr_h)Ѿ�'��C�"�\���C��9�(��a��ǜ��"�@�`�,��]���Iý �<�^��Q�;�ڗş�Xg�{���CF�P��p�m߹C�ҵ�(���k������]Kc��ʇ�l^i�s	�":��O����W�w���>K[ W⃆���$E�<�< Ecȁ�g���̅�i0���I�~�s��f��s_:�L	9����5
 ��v �����s
�)���9b��N�O�g���X2�ǲ1<f�j�5�զ�oUb����q�2L��H���V8�J�!�'{��t�&z�x�{l��j���#,<����md���zWZ�ƶm�öi�-�Js��2���N�ðhO��2@��(�+�n��̄�[̈́T�<��O}JP��d���?}�R@�c�J�pѓ����R�,�қ5OȒ��EVćc`��0����&/?O� }�3oC�l    IDAT|�j�p��a���_��_qf/�<c0&�a�������>5�Y�9+�Ϲ9�p>bi�=��},�x�y�Ґ,­۷�5�$i%�ʧ����߾�䓗�	�����գ[nퟙ<��nX_������Wٖ����A��乯PԐ�a���D&l�N�� ^:�ق�K���t:�@��y0)^���q���| �55�+�eI�</��9�γ�/�Ģ���̢�n��X��n����{���VV��U��5,�N��a5��Z֎�;��!I�j�p�� �e���{F�<�i"��L���DGZ:t�eC�ۤYd5��j;vm��}�c>xh7M"9xfs̩M�,&#�KE1����4�n��IqL(h҇�-�&� +[I�|6'�OZ�9�&r��������=�dԢ���#�����R����ʜV"�/�*�G��:�#s&�~+*�>Ww{� �w�Gڡ|:��=��7֏�p�6�关��q� �w������cz3DNl��E/z�;���	<P;s/$v�`c��"cY�q�ߐF�S�Y>g����_�ӟ��M�L�m�I�r����v�o����G��:�Μ�8�U}+�5�y��+���g�j4Z�P�xb�$�j���x0Y���á�`��������x�
N�����c�G3ؔ%#`�SsLK3��YVi9�ҺmX��.��R�)�Jjq{��{,�����Z6�����*�%V�v:cV���ê�ͨQ������ a_�<��@���C����fU��W�Ht����[{�6c��y�؎];PX,�����^����!:�1x?X �-������\d!���A,	-��_AցE�,��O A��<���m�8�o �v��x���с������~�/H z@�����':��G���x���G?��Ge�2��_���:I@� 7�����d	@�R�3�����I!�$�3Y��8N6�|�o]�d@xŎ��4��#�VWM{���8�t��o����5� ,�S���LQ�w��*i�����/ o�V8��I"a �)���/t3X�k� 7��!��{��k�P���t'-���ε�/��(Z�T2��^�w[4z��'�u&� �V���X;�*@xM͢����aq5�v	��Q�`����펼*���DByP�ØV���Z��K�i����Q�,J|�	�s�T�ik@�I:��B5���̈́+z�@�����2�q�2a`8|��$�[lsR����
��b�k�qA*��s ��b�1�áDԊ<�rl��cɄCfͽu3aƗ�Z�Ҧ��7��1�7n��G;]u�U��}���Xrh ���'���'|&'��QV���NEf���yqέ��Z�ǝ]N�8�6���w^��������j��;o�=�R�#�Fn�x����r��{k��ۿc{��u�T��<�FiHҠ��cN|�;���d^�9A#6��/��l����'��AJ�22�^ �=�q��(`^;����n�;�.-A8F1Ha»-�{��L�rĄYҮX-��c�%�yâZD?��@�9Ⱥ�� �Y+�!�c.+�
��ؒw�5�NV�H�p6�D�]{v;v��qhƲ�	�	��e�jA{����-
c��o��+�`EL�4j�έ��q  YʄY걡�p+�S�E���X�򗐀�sa��_���X�ɯ盭m�N?/9B�7�q� �u�n��O���6,�$0��?�tX+�p�X����q��״��44?���tb�C_@���/��R�7iǟ���w��noodsc�<@���e�{7<�l���n����L1xJ�`Ő�%�=7Xw�q^ד�)�ê"ݏ��Ӈ?�Y�t�M�'�h�l�'g _��>�B�T�%B��l(����S�f�����B��jn��a�#��,۽���أ#`�E%Nz� Ѱ
L8M]�)4�"Y�x�Cj0����d�I9��������׃ӡg�4 l5��9��>�яt������t>��оfa�c�	˯�s�Q��I$����d�md<���BR	��c	�|� J���XwH�[�O?��uc*S����Eb���ǚ	�ϸ�L������w�	kH�j�P��i+B\�z/�g�+	��"��t/�"p�9VQ"�M�0�JQRT9�r��]{���}��q��y���Q���P�jN3���U���/�c��ۻw�'+��t`~j��0����d��<���48C� F������Tx	�F�����A<���`Z��c��#�~~5�ن��y(�9@8j�#��{��=�-3���,A����6c+V�XқZ�Z�	�{Z2�C�ps����,f�T�פ��4�Y#^i{��>��Ԧ��1%�k�}���T�͹Js1a@9��	?� ̽�AĠ'.���������cG�C��c`���`�9�T��}|��G�3�I8�]8� a�5!�<�����_�LD%�������!��� bƳkLз|/Y� #sN�j�n k�L�B!���q"|�aI�\�q���u�D��Dj���y�F�����~k�Ax՞�n�Z�o�Y�*_�o�y��G�e�\nO}��;&<������(�a�_q�����XB�-��D�������;5�u�D�|�΄��S��>�U�2�(����b� �ǹE0�ֈ�,Ax`�f��[2n�kWc���ZeƆ��&��N����v�.�o=羞�QTS#"���URSw	WJM�hOk�LM��Շ>��t�9��҄CGR8�5��ßgt����,�)�i�L�C,1$
�0�1@VĠ���9� 	�Ysį��x.2�p��_p����/�Y]�7>X�9�[��$k��m�I{i�S,�p�=�UD6�X�)�X�)�_�D�(� ���H��e�b���gL%I�믿�ͧ�vZ�f��W.B���?3���6��!k����#���ϿЫ�T�&	Ńk�X�y`�[<�8�4�@�QQvV:�A�7�/`��8��C�r����}��sˑ����9b�q�!e0W�#.��b7�Jdyk�V$;�2r��>`�.�plQV�V%����:m+�L�A&L�Kg�D�)mY@[�����F%6�䊈	��	Q��m$:ڲAs'�t6XD]X�Μ}�`�s9$�c�b����v�-Ą�cN��B��h�D_�rR�����B�L=͇n=u!Ki��h���}bZ�З��u2��C�gZ$�Gat�Ƶȅ���d�z���&|�SV��WI�q��9a���r��>�`҄2L� Ua�*����5�/�o��^K�\ߛ$��������SNپ�q� ÄZS�Z�EloT�F���N��Xjδl��՝���Nx34�J#�aa-���.�ք'U�X��Z�X͘��A�j*�.!}�L8�T-w/<�#S�p�:���+<�"�T��{lE���?���,ߵ�*�5/{�&�5r�iZ�cվ��6eq�>w��Җ�+�sA��je��q\��OY��cʆlĞb6|���������d������G?�1DZ�d��jr�=4i�R���sK�q:<<f���Xf�&�)m��	� e*�1�m�p�R3��g�1ǘ����l8)�pqYʄY�cgc�ZS��-+�]�q��r̅���sR>�;��?m���e�"�[9k�gQ�V���\EbѶS�1�P{�f��o�qE��0[,&$Q�^�B �(�`�~`A��$�Y��9�ƊA��P�?n�⁤�J4g���r6h@i i ���x脜�/%L$��#�4�(���iIԴ���%�\ayT�(�ytĊ������F�|�KƫV�H�Ȭ�p�C�*}��(�S�"G[^��K[�E�(k\�#��&Q$8Sʒz*�3���3,>�Z}'8[Y�~ddrY@�I���c�Q�θO0 ���zʹ�@�u�j�Q	a�j�j�9M�p⨏%K�\_s,�� ����{����\�x�ɿ\�/'��_��x
�R���n܇�Q���e���A���b�b�ݖ ��/�
#���f9ڰ���-�p��И�Y��H��2�3����2���~�-��/��/����u�-���	�\c�2�wZI�h�������Ԑ���JիÀT!l��,J�Q�7��}V�����l�����c@���V&�,��c�}�l�N�Ɖ����0��,A�m�h�ab�Ҕyw��>\�1��uΫ�!�"��|���3,[>ѦmЬҶ<�ld�1a&��61dEcU�"\h{+����<�ؔ���K�FAh:s]9ESE�/���1�!�-3�X�/��J�S,5��D���̧��a�@�9����zDu&�8�� _��cT֡p!|v���/��4~��y�RP}�ꫯ~���)���d����<�4�pjUY�����%J�����>���2�H9v� lYW-&D-�a�L���"D-�A��ȧ-�4l�0�p� Wr��,�Ȏ+�E˨A�����Sт���F�ϩ���^{�e+N�f߉6� �~��ޑ�b¬����M�y'����j cn�?Ŵ���9� �|���2���=F�_�R�Z��.�*G�sD ��e��|�X��
L����+��\[	�}��jĜ�[���	/�8�!�MC��M��h,�3�|�mY�a�yI��tssi�����v����F�đ�NTCΦ	k%�3��.�@���>$I�˄�j�~h"9� �K/�ܓ!�J��ֈ��wX4r������[gUK) ��XTi� L�ܴ���R@�eׅzV�q&iCr��QA�cW\`�$ =Ͳ�S����0���yj���oM&�IF�$t2���>X�ژ��!kcV�_&��JJç_ m�C%� F�T(1i��g��Q�D���	/��1�YHHr^��#Nrڗ>�?#�x����A����1"���>d���"�K�-/dg;&���tȴ�H�� �CK�G�<z-(:����&_z�;����g���W"��	��6�&�Tc���� �!�sp���39��%GT]�hg0��ˊ�JdI9b�%#�Z������'2KҚeq�Y�� �#T�_���˗6��w6�$�W�k�gЩ��d���FO�lų��m� �,�ѽ{��f���^�2�F�T{j�G���)9�|E�p����`�&6!�h� �����7�^�0a?���>Iԑ�|���x�\�+���0a�@E�f tZ�	i�(���8"p��
�|���x��F��6n�ܦϥ�ӧH�:Sd��R���$-��]J_���l�fr�"fb�]-�"�)ZV[qLX$ܢMU0���f�{m�j?�Q��kU	�y��р�*�P�;�,11�Q���B :"�+%gv��뼞0�I%�>+���z��l�6�ɖUҊ��m�M�jᘫ�1iqMv[TM+��[��Ow�#.�Kf�;YSLq�&�a�c,_y������h��fY��Q@���̈́e�2Y����U���r�i��M�|���5�b�3i�Ì�WIH Oz��)r  `X8p�!�(*JYv;�y��(�N��@����!X`�B`����I�� QO�0���F3>�Ѩ���o�)���`GG,��"',V�~�n��cDFĞ�\Z��`�>�/_}�տ�sg��u5��թ[��i���!u�:�������D���`��SO��CmR�G�����.����]���c[,ݽ�l��!jq^5j-��=V#m9���kl Zh�*a��j�o���L�D̡^���m��\0e���h�'Z��X���Q�3��>����4X%�҃Bט�r|Jv�x&.Z;(8^+�ˎXv�Ez�yU��3R���1�n���:Ąa�%bQdn E��`� ���N�d�J^�| Y���IW�{J�R�������S���g���.�Wu;5�ĈC|���*`�v�q^����C��F�`�c���}q�u�V��&�LZ�S����aM g�e�p]S��YAè�j���|v ���m|z�*=��f�%qfg�;�֟��B���6PkXOk���wZ��Vk�|��vj=l5?M��*=��V�ޟ[�PԽ�l7.����
�}#ϝ+I�>���~��UkE+m�~���Zk՟b�jeв��G?���zM��[�_��~�U\���M:Ҡ�6���H�..���Ċò��$�����������c.�ﰟ�]
�׸�<~��)r!F�x�<dRr|jQ�I;�a����J7�}��-����B������=Q1�$%-���{~�%�cMDI�����g�kt��>�YdOq3ܛ�l�w�Eڂ�BB�=��Ӓ��x�oX�d���4Ԟq���nMb���g�S@��0Uוϙ�ܸ�e���A\#��al����X�a����^22'.��g�L����f$��@�������ZW�hU��b��"�!�	�[���ZwHXk�U�j���T��ֺ#n,!�(��v��������͏;s���0A�>�<�ν����y��|��}�{�ѓ�jé6<���+͟�gޞW���J�f�ғ?2�������4t�})�R����fͭ��Y�)U�2���Ŏ��O��;͍.a.�p��G�s�A�[ޏTSo�i`d��뻺ӷ~�5���z�>4+oo�?0��fW�wݞ��pΧn�b�A����ٌ�Dd��@ϧ�R����ar �5�/R>s@ǙT�d��B:K�C����&N��O�y�:���s1�`��1�J�@X������0�H��m� `��;֔���˾k�5LG]���0<�L<rue�jo
ޭ�8+�3 �A9�� |�����-����h���8k�O�B5�.� ��wDo
���W�s�_5�5���R�|�Bc5>!����T��I��q@`7�����Cs����ݝ���Ҳ�H�<|ߔ�ߛ��G<YB�!
����9]����b1Fa T�h��l�+q��k:X�\�J��4R�3m������Mw����4�wn���<��I�Q�� ����YC9n2�e����HhG���mTpqq�!m�̲��g2cLؕN���;qO����xV�F�q5�u,�8(f[��j��X����`A�v�(Q�6����x�5�hg�qħRg���{%�8��?JأP�K��w�H'���1w����Q&��'�y3�ޡ	+�\\P�a�N/bt�9�����gܪ�q����1A8�Sȫt��z-k��*}i�V�	�{�7�=u�t�K�z��<�r��Й�׺rv}v���~�#�d�����0[�0.rDd�ݨî��H��oY�(r���M��J��3+�5��`eϼ�ܬ��42ܕzq*��	��;��ul;D`G������y���'׍S:�����ц�e9��x�x?l�)5�F�|����e;D�}�m�q��� %��I�siyd��c�D;����+��}G ��y����Ĉ�v�s��&��vm��x���0ʛ�m0JL>�q���:����3����4ox�ɀ0�0;k�	Ä��p�O;�y���J��p1���r�Ƒ�ϲ G%��wݑۥ�+˶L� ~��s�B��,Fm���C�eO�>�����Z���	*Sw_ޝch�Z=/ި�i��)'ú&\�z�����	�yϏTEbIi`h0�V� y,�����ޑ�T�w��=�RmhG�&�N=�p��:C��� ,��ь�6|Ɏ�%�C���dJ���#(	XN!a�q#˩v��:_)I���"HH$�t:j�x#��b�`Tn�g@��8˱�c[ęQ��9�_���t�o�{�A][�;,'��4ͥr���qF�����ׯ?���,:�m݂&��2תEn�rr ��I��ȍ��J�NI�C�C��	�����F�GϽz�w�0�#�E��0�X�Z-��HwW��3�D���ONVv�����W��9�C��v�V�'��x+���H�N��ùJ��m    IDAT�r�E<p��Q�w�``뮧
@?RO}LS=�{G�}��4������ԗ�#�4<8��K}�l4�8��٥��LB���k�Q�ߨ;�3؟�E��i���kp�ZN�}6ʍ�ow��S5`m[���R81,�6�2M���(�U������	�n�1��o,�1�Y�`�-r�a�ܡ�R�Xvن<�P4%1��` g{5�0�I��� �c �V�����	FA���W�[����a��{��-7]6���ı@�o�G�$��RHC������O������
�����n�ǘ{�D�q�T5=�c�
��@h �f�uో\�Y�������Z����,��\�I�������`���2-'>���`��]����袌"�ew���ݬLN�Yը���]i�p�W�){�9���T�	�y9��3E�����4_s��؉4���O4����S:�:8���I|ﾲAX��Fg4�Eu�������v1����m�]��x Xx%)�7�x�V�C���f�Q��Ⱥc�&[�c1me�Y6:g�D��O����a N�û��㽭�Z�FR�O�]����not�)o|̂[}ټၣ��#�,MG�<O{`�,�t)0@L�#��,����H����F� ك�կ~uf�9²��_�%}����F�lC��:t\l0�����@�DO7aa���RO_5m��K�>��ޮB��W
�2�YlW^��f��sNI9�0����bۣ"�;�,3Lf�gw�kp�t���*��ix`8�)���]��h��3Ə�k QFh�c�'W�;DD�O��9U�N�DԣǺo�X˯3���d��8/- ���h)A"z�%b���l���9^�ԁz,`�H}4c�9?ړ��l��J�2�";��C`x�@\߈+���X2L���$�'F]���稍�GA�̎���3�}�­7_6����f���������@魥�G��z���ܹ{��}�ĎJ�!���cB� 8a���I@dtTSw�[������8 ����,6d�Ҙ��[��e 娅��JA���ʷ��b��w(ݦ ���FW�!d�P���G&��.'|gq�+��n�1�sfj`���8#V��oH��t�Ȍ�-��/�F8P�q�gnԈ� �0Y��y����q222R�V�W�^����������qo��eF�����>�ꛛ����%��}.�g�����<3Z ��;zEu鄃�`h2 7	?H�c�Q�6��F$������Pl�Ɉ��h��2��t|���f6S������j@)�߉�!18@�~&���0�S��3���v�Q��0��7�*gI�3GI$��N�Wv�t�pT��U��O�Y��� |���{���n�t�T[>8ԟ*�=iN����כ�?���'<6���?L7�pS~xG&
�X�W��2��T�ёyg��I�u��(lEr�gf����hv��yի^�+��@�0vT<��L�����=k �����/��>�����ӟ�tƒ�N;-�ڏ}�c�8i��'P�p�	YZ��%��o����p���*P�o�t_&<��U*��֬Y���2a@x��o�t��m˙2�T����ZZ�|Yz����n�rC����#�2Y�:#�9�@N [�8!��lO�6��xE��9�5�C�1B>�y��K:/���V��{�}��5S�����V5 ��߮]�6˖��H(Dn����gdݖ���o�L\b��g>��!���Ȑ�W�z��椁�q-�y3 PwvF�X�j���޹��9��d�	���+_yR���M_��������<t�=��fu9�0�0
�;R@�'��e:�ta� ����f$#/8�{���8H��V=��L����Y�k�o�ƍ9���?������s�T�d��ߌp@�$�j�9���~��8j���c�0��Db!��?��$����3�Wz���z}���s�ʋ.:�裏�c"�9��Fh���vå��+�g����:��?O��vk���'��0� -q�)����lt_""m[��]ՠ��b�w[#7�|]2��f�੠�,6.��d��D*v�ؙ����� }��~�Yge�ǌ�+_�J��t�Iy{�ؗ�����~p�햸; �n�`~#���J S@��	�u$�Fd�w�'�
}�=ц��ow1�p��犕o��G�a^t+ <�"�k�w�#Z�^�����~�����s�c3� � �a6�y�o��%nh��~�s�˕�s���>7ꄓ2�u�ע!�hB��͵�1�i�0s������	�N=���p�%�4��������H� "���,�e��A3k�M+k"}�S�p�br� �W\qE�>�ឞ��^|�9aC�fo�gEo_5uwU�҃O/|����?��t�/�z�}�
�ٳ�l�~�2@�QG����k�"F/�7�q%
�d���'���m�љy��)���vr/�s��㙹�L����k��f��0�8q�� ��_�H ]�3��
p� +�~�QGe�fd�=@��dʞK@ 8�}�o����+�+֯[wnGW̱Xc��o�l������R�қ���)�9�yv���+;���B~ (M�e��Z����<������+���Y��-�tR��Db�Y0�py'ͭ����L�&w��؀+4[�4�+O�r �剋����&w���fj`�5�bR'���$�����~&h��)�a�G� 4Y��~����Z��֍�pI7�s�x��g~��[2^�j���+6���Yf��n�l~}��=��'�bɲt�q�������0�,a m�/�1!F�&L��f5���e�\�E�`ʡW�� Yco���Lu�Nfq��IE�+��d���yqE���������@���g����]Q�#��������P15Z�hq��C� +�lGb{��h����a���+s_��/��8�8�.�i�;�w�i��V*�׬^s^g�#N;瀇ܺu��{�Ȋ���i�cN'��������?�M{Ι�����a��v|+���n�v������O~2��6c�,��F$e�mres'�s��
�h���I���,Nڽ�T����u�KY16�nq��<�{Ϝ;SS���J,0��MDF�Y��=&�r��/� 4�4\���0�p�o�;���D]�w�e��&������^A�V�t_�f՚s:
¤�|ح[7Ww�Є�ki���N:���Gw��7�=�Tzs�'t���&Y�s#���k|!�Þ��?�3�ۿ�[�B ��s��:(k8� F�1`׀.e� e�;�	�G��Bx>���j��:�����['N��aДGО�#vU��\�� ��^t�EY����?�#�d����?���o0�Q b��׾6�� ��nr�{��9���H$Տ�vf��)��ȘE��QЮuww]�~��7tT&����o��{��O�ф�Y��c��yp����t�w���"��K��� OY+� A��d��J�2�&¡�4�!`�nXhs�4䪫�ʂ��J���54f hW��PN��N��v���� >S�������������vjv�]Y0^�[VŲ�����l�1c�g�}v�	�����Fg�`;��&�� ��A	��s b���I�93(�b�.�Q��bnÆgw4�;�Ϳ��s��S�v�sC���_�����$n^�|���
Q(u�Ȯ���p<������ׄ�?�ъQ��/̕�bt^� �ד��f�\	CÙpyW3�VH���it��1���u&�{̲�5�z�_��;`\^54�	O��g��d�G 
o�۳�K�6������R�>��<�Ɩe�XDz��$n �a����q�]�'�;,��C̈́�%��G��q���wt{�%����o�_�JN-�F�J�?���)G�'�����~�n�qK�XP��S��0.� ��̱_#�3� \��9DE�(X�3�1�?'��	9do�����a��"G��-o,�I�mv���D��`���@t�KYC��e���L�`�Vlذ!K���Ӻ�;F��ۿ���س)���! ( 6�G��G紤���lj�#G
������>s����y��כ�=�,jh��g�K۶ݗ�~��t�I/O{�~��~��F!e�N	F�_�# ��K:K����_�r��-�y�a�/x�r���5k�Ne��LN<��� �o�FFD0�.ӦL�>��g���ەe�i�d�Tˍ ����͙����Uf��n(��L]���`R&'��7~��,`��'V�� 1��b�[臨�p.�{ Q��#����(�����ի�\�b��v����]�����7e9��-��3��N��f��K�����G�I}�~���0��.tH�V�e)!���qn�"�������z0Ss
��%q�X 6���#x�r:$y~�ɑ�ӌ�q0������kT��1F�-����5���
����=^Wϲﭞo"���xl9,��R��~��(�Y�гo䑳��F���{�R �v1f<ΞʳJ�#H��m�M"��%쬁4qd�da��^�)���8��� *)FGv�Z�z�ʕ� ��nټ��}�u�����#��?-YrDη�*5m5��Ί
�~K�(}�m7�V��^���F�wݷ��T������Z���t�TA�rǎZ�.Q'�Af���!vJG�<��&�',؄�+!ŭ���k��xJ����ࢮ6è[[����8��Ȩ_��ٞv����a�!�dL��nx�mI��6NV�QB�OJ�F�����$���	[X� ��.���?���!��f�h�h��F��.ᅷlټ���c���]��7¦��4��������ex yHqTعy�^m�(�Ȥb��=���P1�Л�q�2Io�6IT6��ow0���pd�J�*x���A�E0��z.l��L�S��1F��-��'	S:;*���L$�re3Ze�����|Yg?��>��ːe_q`��9 ��Vl�����,��
�'���q�v�ߝ��g��]�������h6�C��|����E��o��	Q[x�-���C*���Hv�U*�y{��jW�>��R��E?!�������Kv+iTP��9��ў�q�^+�����Kc廨�L��L�}��F�)�O��m_|n;��c,c�0{����k�S+CZ�aꋲ.�tNɇ6a��3Jmۖ���3r��V'����2U�Ҏ_f��]<�w#����A�ߔ�l/�]�����S��о֭����)H&�G��ܡ3�BWRg{Q�Q��l>�jժ3:�	��޼i�4�CԈ���P��+�y�{k�l���
��x��70�w
^��G�|���]��q^�{E��4��=;�Qv�^\�5c�.q�ȭC�7"�����ĥ�tv��#�N�G:A�rQkC�f���#{��Ap:۾�{��r�38I����?���U�5/�}N-Y�ٶ�ɸ��rRԊ��(��ygJ�_�g��c�?S�֫�R��D2��,�D$���J��yΎ��[6�ڞ�p��I�ၴ=��k��OIc�Ԝ�8*;hQ�N�Ai�\S/��0��זEG`�#�*ǎ�N�@�B.�� �p3:��Og�dY�I&�(�jL��п�y������~G��҉��`��N�M�{J:t�Z��$5��Q7XW��������՚�f5�2�*)	��a����˱�M��Hg�;�	��y�������@x��n!w�15�UO��	���L8�q����O�n��4����5Em3o��:�h���ָ��8�
�ց�6�8pJ���{ �a��>��G��� ��.f�����	�'L ��� z���Q����v�{�ʜ�҇�oY�ˀ mI�	��� Sf�T�s��>��������Y�ǎ\�GR�wfBq�Jh)�%�ҁywg0�팜:�e�\g�b�����,������R���U�N�a�ڞ�ێ��Ɏ9�-��	�h��6,&��,I#��� !�Ƒ:N)��N:�1�?Fi����S��`t*HG"� ̋�ynS|�8�!lQ9��Y6��g=+k��I%�&uFAX=��pʱ��N$�)��κ0�[��e�W2 J���?=�����G�đJh&Z%[��,D`�5�g�����Z��c���S��T��0��ݩ#R�������X��uhc���|NyIሳJIbw�g�$1���sٯ��R������Z�~n�ʕ���7�ߐ#p�EM�|�lo4�+�k��>t�si�udgN�v�!��=Ǻ� [�3Q$n���;K��q�-��]�/����A\ո(&L�PLØ�u �h�>#I���eS�9"o�z�U�]7��8c�{�'rvz���������%3b��SN������75�K�_���e��o~s[^d#�"	�7� 6��~X��C�^p���X*�c�2��h��I'�@rg��g<�`Vf���vlD"!��>�6���[��OG��U0�@�ddƞ�3�,����V�^=} �(:�*v�8-K�h�3���\�� 0�����j����@
`	[24�����v��rm3�3	�x)FX��&d��> �&�S�k�0a�2jSiߩ���p~��|֡e��$a�h��?;ǰ��$A9L�A�#�Hc� [����`�.�k�\���xΣ=a��S�^�}h{ڗ�|�0�^�r�=ǐ��킢��l�ϱQ,��V}��~����ҁA����l6bV�Si�f��e����իW�:mL��
��-m���:[�L8���P��u���a�9�IX���z0 ������d(LU�6�9:*�ҹC;q䍨r�B�AnP^���7\[�w=�s�<e��� S��v����ߣגf�J��A� I�=�i���h����m~Е9����r-]~�3�%�����n�àMx"�Jy�=8�<����L���9���� 2�2�;x5g�o����,"�h�e�Fn�Kwww�A8�	�~��yC�O6:b,9����� qA�U#8����\!��P�*6B+&���Q^�̹���	�+�|yǠ	�1 c��YB�Ш�{����q a�q�kP�g̯@�W]	�DD����Sov���:�6�kE���I=�qw���EG��Xe���}۔��3 /�~�����3�5ϋ���V��
�9β웂0ύ�20�~?Q�PD[�n� �#����s<�Y�/�p3v@��rI�m�i���O���'�v�~q����oy ���*�,NכU\������@/w�����l��tZ-/?�n���~�ba6����Ɂ�@�5�N���AE9�c����܁t��=\�)@������O[I��TR��xw� �m���$�h�q���b���؆�q���oAK-U�Zߋ�t�ǁA��;�C��bߚ.K��-Gr6D��3;�)Y��r��>��������_|�i΢v����qæy��O���}F�q��fc5c�>���]��@��)_�ȷ*�n��ǁ��bGta�L��b4�XSFt?e@�Fa���D��q�n>˰"s��щ��g;gy���;�d������:���d�N�e�����`���]�F=��D�1��vv�qê<��8+⻸�7��LT0���#���a����P�Ѫ��V<>2kYh�-b��e��s�7�'~�Z�Hi�	��&|�ƍO�hRw6�\��f����@��M.�"D��м�HV���)T��+O#�M��݊I�j��{3@m��~�!�r5�������}���L�-�h�YM����0��b�ttbK��[Z�N�k��5T�G�=ֽ�S
�D@�H;�>�0m�2X�����]��\�/PF����w�j�\י�������ϙ��Ug0�%�����=Nn�k    IDAT�˃4��Y��"�Ł���@O=(��V��2�6�y�#&�Z�8j�J{�E$�M@x�T�6l8�� ���s�ϖ-�������Ã�T��Ô AB��s��E��e�cQ}��Z� ���S�����"��G��x�؋����	s0ؘ��%�t^�&E=��3�Y����&�-���=��*I����M�������E0�Q3L����zR���U�V�߸�	��d�q���UG�{��j��G�$c4���pu`y/��t�U@�r�dAXP4N�ε]`�w���l�W�tf�5�_�ڙE���c�g� Bd��PgQV��������������s���?��-�����"�����ܞ=ROO5�n���7�7!G,\�o"'3��놝�)5H2e2��a���9u4�3��!5 8�xVxq/��˼;��G��`�>\d���
�W����FA"{�f�jO��k45�hxh��>u�P��������G�Y�L�����APo0Z��9c���(/�e�갲R�h���9�&S�>���;�G�)�DBP�=p�	^���:�̤�}�M#A��z��.3β�j{�g���@}�x�xԩ9���I��a��=���l�H*��%: Z�>��o;]s�5��2(��� B�����3��DT8�44���^,V©N��"���y�Z�>
�gv�;���������I�#��R��''�a�2��k#�i����'=�������
��蘌^T&�H��*/=�N��n�R��SO͙�	��J��\���.��q=;�#����jw�N���-�>RhIN�uVݷ� AxpT
�1ֆ��p����k��f�ޣu@i���Z�:.ue�.��Da��brωr��Q��q��q��u1­�b�AX-���]���h�/�}��
^��"(:+��	�Ԗ������@��B����#N��lZ���S�X'�����@�5V�Z��г��5�yM^<"	S�i��#yP���0K��4��[���wY��XZ��KRJ$�v���C�$�[B������n�|����f�\��g�s�q�\Cs�[jw�"4����?�fAt���gW<iߘvqϬE&��<��('��Â4���"B�Y��#o�02Ȕ|.='�(��]5�I��J��n�E+Р�˿� �IK	E����!E���s]ų\�&�}Gu��q��|W�6��a���;��&�Wgk���=��C��S�B2����燫�U��+���t���SdZV`�l�O�}���$E;߯�SA�A!�gGi���f^��G�AEY]B�8���w�Z����6���;V���@����pҧ��ȭE=Iۍ��;d�1���	\�E
o������.��]_��ɾT���᯻x^��ԽO��@�1��<�n�����xĥ�D��k�ߴ6+���,���@�a�8��7�4Qf[��|~x�J�2���e �4�g��ѩ�]g[Z����K܅��C�A��W���'[�� \e��@��G��r?Ti��~�D�;[�ǆ�|�̻��	�!�L��m<���P,�ǈt⺪u�_t�D|�d�>���[M���@g`;�/U�:���6�zs������z�r#K���cq(���`p5jG[�
HJTS����b�z�$%��-4��6t��J�������#�m���
������B��5�C!��A���2-D�V	��/��߯q�0Wo7*"����?r�oi|��x0l�����v+g����gd�0�E5.�(�U�Y��6A�z���卣��pBq�[�eF4Q�Kv[Un�D8�;T �����,�X Ti!�#HZ�&,�K�<�u0J"���K�� c�v�!����y��!E��W�m��|5mA�𝌸Z]}ʺ*1~b Q��	�Sv�]�F%�Ҩ4���/�q ��R�8
��Al�M�#�7a���0�Ã�ɑ�>�+~���~�0�����������9���i�<dF|�)c��R���f����s��q���G$־�ݙD%!I�l�or�&b��i-9��D��?�{����I8]�����h�&�H?������ 4c��~��j`壬����+Yݴ��z�lL	8|�SLT��}�'���H��������9|V����鳯L�! ��{��������Mϡ`
*�e��V$8�O7�=�g=3W;���Q�M���3��o�R�,�>p�;�xS*��g�^�j�g?���ѹϰ�0�ik���O��p����]��f�V�ǃU��'sD���{�=����Ue�±���-�2{�^H��� ۆo[���m�����+�_��EAA^�U
�����!(ĿBӯF@^��?*��紉�P��:)��/�� ~����n���N����öQ�*�H�_F��}��!,���bw��Wۖy��}deQ��\C�`h��(���+���_l�N8w�Sد��E�6��%�6�e�§#���_K��R�v�O|��Or�?���7�-�a�*�z<GĹ |�BL3��D���c[��0�u��#�������!2��J�G{\\\GYY�ί�.�
T>}�lE�F�Iʷ?�M�N�o������$���ةA��E�f;��L)Y�O�a9�6}w�,��on#�\�P���;P���x�����/�u;O��ZC}�&�~�������;ym=YHZU@
��y���NOG���2: ���̴}�v�6��7���"d�(#���h�&Z0)�X�_��v|؄�N���|q0�T�P���A'`��0z_Sɻ�X���C�f�m�����
Y븀<��̠n���t%�	���d�A���)/ e
�US��������nMYz��v���Zf�D���s �*p܆�n��]�N��p<��� �����]�Y16�OpQ���.OIl�sM����п=7R����g�iv.�o����}b�gr��M����>��C�i�mq��6�: "�ɢM�jVH��,�}&�f�H��	U���q�]-���͉��70s8�%�dq�+ű�j�XY�x/��5m��;�����8���������?��B�ѝأ�yI����"�m�y�r{G{�?A��N��}��^3eR��"q�(t���?hP�U��a�&Q#3Ħ���E�nN�x��'v�&U�۬#W�Ϧ�\o�sa(�k�Gh�O�T�QWS2�Eb�zB��c#��$C/����(�v=v=9���u�Z1���G�Znj�G\�Yp΁��wT��U�H���:�#�BP̟����C�D�����u�׿v9���F��G�U x���HV���j\WM��a�-��G�I��Ԙ��-m��/m���UP0v�,z��>a^��Ⱦ�z?ز��S��e��Ci�ĜK�4p%]�N!�d�Ϩ�BW ��k�����(_�V3G܄)��5�Yj���!�b|"ѳ#���UTTދ1��r��2��kP��N�i޾�$�I��^�A좰�.rf��`��8i�*!0�y�?X|q��6�IɲV3��{��O�������y���x�Y%���=����FoZd?K�~��
�����C�����{A~+���5ӂRw�ٸ*�F�o4�7'�{ �{�N���Y����O�4D�^��c�y���"�Ju9%W��ra)��]2���z�!��D��Я0���<�x-�ݷ
�3zܐ|����Wh�x��\����D���J��AyEx�1@�(�q�c�1�C�[!V OK �C���*����P��И���z�� >.�ht��R���%^�@ no >LE%��d��wx��<�)N�y�04>®�|q..E�I*6`�����(�Z��^k����w:�Yج�o���KF��-���GP�X�uM�c����39@b�����=��� ~M��G3�l�?�
JX����"��5��ʡ�w�vC�&!�2��Yu�����wһ���j�ޥMoy�/�� O*J��ts�x^���(l�������k���.��������Z�ގ���M�%4�3�p�+����c����}��8�����µ������l�q����Y#�z�X�������T6��1S�������g^�u��j״�a�_i2�5&Ry b8�?���i���QLݡqn	D�/mZ&�3eS�zJ������;7�<x�N4�Bj�b�w����|
`�Y򐆈~�!T{�i��{��]D��.ɼɹ�zZ+���!�"aJfQ�}��/Gc�lAP����Fc��%���y�ڀ�����ii��l�7���SE��;T��Z��N��p_ޟC����x�hg���J��m٥�;�qr�R��e-%���xO�Y17"h\�F&����:�.yT�?���Я-�K�S��'�7��
 PQ����#�Ty�9���5PJ(� �TF�����F{p���x���M�[D37~�i&��'��Mrnʫ�v��B��7I��c�ޒ���_����j��j��F����}1�`�x�'�v8W>��j���2F�?
����
FR���h;bo3ڀ ���wjh�m@�yS��qV�k�;��2�m��1���W1�p�����7�����8�K�۴���&�O6�/��h�f�����<����}Np��N�yh���9~7
y�nM��.��K4�Cc��_F��Å;���(*m�^|�}���2��;A>Ç�,�t�a�s�WD�EB<�� $�(��^c2lyD��5�U�5��fW y���"�quޯ�+s<���A/W��֝��3ٔ�5���p��Ev�ߌ�^�TD�-&=��+%"�k..�Q{/��B�� .	���"��˰�D�һ5�W�1��Bbn��u���{X���rD��o$�t64I
�pV
5��ж���Ñb�
�_��'}�vd_��2��|<S�Bg��>�HV#���4�v"s2�g}�xu���Q�,;+�<5X����ż-2�* �jܒ�Xy�zff�v�v.B�>��3Z�}o{���*��8�z���eі��ڙ՗[��8�h��	@�@� ЙI]]�!�����A�g޽�c��#����#����z���VBՒ��]h�n��//��	>7�+(w6���ƣACcu$'=j��V0����&��'Q��)��"��6��0XP����D{��ǤrQ���QX��n��g����e�{%`?<+E�	������ID.+D�,d���պ�TF�^L~�^~�A��^�#�^=ZV�	O��pS�=j�DF���-�1X�H�I����#�W��PS1�����z��.��a�a]u�h�@���;i�.P�<Rx�>c�<rr���19EGu�l��X:Q�d���� ��'�Z��t�g��'1��?.T<��X�V��T&&�2�t����?W��kȬ܈�K�n�S�;y��>N�%��R�N�[�eL&�|�H�O���{�t�D�h��H��wyZ�6���T�)l8e�ǭ�v�ʂA|�&���Do@0�juʠhI�y}fja� G��a_@��^��Q�����M����E&}R��T��7�,L�pS����l�c}r+u�r�{�{�]�5������(.�&�ޯ�	�M`<f����A���Z����~{c�������	"'ᬳ}���67���L��g��ɋ�ɩ���%��Q֝�&;/��eb�m͎���ެ�WZ�5��?�7���|y����HFF ���>�Nm7μ�a�`z|GB�J��v��7�$3-�i�����m�4!�2��\�O��x� Aq�J�m��$ͻ"��+��f|'�u�
�6QH#j�r�QM>jV�m� �<f�b�w~.e�ёލ �j��*�5-.g�1��ss\:�3�+O�|����!L��K?�m��
��毉��׮1�q4_/�1
	�&���yN�,�%C�F#/b��;�b�`��X����I���֣���0SK�b6�p��a��0�8�/����w~��wL�y��5�Rgo��^^�(ѹ���:��I�[@��Ո�a�[�I�ZӨ������j*�|/��x�\�+׺^O�雏'���dф��ao�^� ��T۽%��An�������oS]�el���}����~9�s�f����!�F5t|x�RI��L�F��O%c(`��A�O��|:\ɸH���7�&�X�z5�R�di�$��>�6j�������s��A�$ه�J�{������1�<�N���O��2�J��Z�6u��񱝟׉�OA9��Z�����|��lط3S�(��ӲK�NMem�ƅG ���=�jX|�URr�r8�"�&K��\oU���XU�O!���u��(~p�PH�|V���T�s�ƚ?>����A�)w#����nԭ5����LW���z0�0�"�8{X!~35�����~"%��ӕZbU��.��3���eKC�Ro��/s�i��zA��j�]?�Z�� %eX&�b�
�֗�����8�6l��J��� %��R31a��֞�N���IT`��]��Ĭ�H��W�j�2�V���n�h+�.���7)�ғ!�3���4AT����&.�7��9����~�װ�Y��ʢ���ќ�Ƥ�B�,ee��@lWHj��mE�	��G��3�.���\��EG�'�w�o9-�0��s��{Z[��C�jh�w���K����S�>��an���3��o�o� �fW�^�	��d�V����R���<��P�C'S�߇B�lBV�p�� �:֗���V%or���mݥ9�]�h�y��2�G]qndBs��L�FO�p�G"*���5ǝ����M-��W�|S������\�'�u�BQ���t��8���pu���˽&S����q&5�v�����Y�]�'��Є�w�ʒ��l�L�Ge�S�����m ���[$�K1��X�Vu�ϖ�Q2�R�g�F�ކC�ّ���_> x�Y�p��ͽO����ș_���fLUhfH;V#I��[1�(���IM��˽��B���*��C����߄z�� 4D�葳���q��]G����z�;�'���.ݼ���ⰰ�HT ,M���`����O�f�V�寍h�6^A����(���t+2h�b
�"����_�!�h�JYx��W�ϵNyo�C�nu��>B,ۤ6,~;t`?���]����M@M]P���"x��ۯʏ�� t���T�o�P���3�����掟��0�1���tK�[�۶�Yr��D�~-B�&�T�%�u�k����l���IO�VA��6T��:H��	�?l�$x+Ov���e�S����g.Mt�3��K`ͥ��J�/�4�N��}0�{S��n�/��YR����� ��^���@��7y'��Q�T!��o���HU���3}A��d���y��K&�l�/��s�������5w@�[i���~�A��� ��,�3݄���	�6�f�M��ק�X<��m���~�~��X0J�{3�D�|� t��H�������)e����P��H?��O�$���g�>��o�oa��s���I���h��#��|��v�)1�,������;c~�Yj��}b�N���vK3��0�O[?��l,�v�T�|�sy�x���G"7�5)X�O��jf*W�y���ﭫ�.������t�Aliҭ+�&j)��1NB��((��=q=��nR�ɦI���2�rȲ��j&����I߸2gc	���������H�y4bY9�����(��w�˾�t��j���;�k�`dx+���{M�JT�������Z�l�t���|��t��\��&��}�i,w3]�c+��?l%���m�b���9g?%Yv������LV�Z�HϬ�^	d��������j�J��k��x]�E�n�X�E&6c������DRZ�i�B��S5���ug��Z��'h�NN�0����4$����\.�{ށb�i���h��
�Y�2��Wr6뎥$��M�0�7"Z��Rs4� ��Z���O�88%�ʫ:�����4� �g�g#-��ڎrӳܾn�Bax�iȷ����`H���ϓ��b��׷�7�J"+/0�O���N���AQ5j-�ž4��y��xQ	���$)��.�?�b<�2$�>a[g�s�����_��:���zZ+�8��g~k+�X!�*�_;��\������	�B/ �&��ө"���ZۂGנk�0��ڦ�_�KSM�`�>�n\�A$�mH��.�ؗO�C#.�AQ��Y��ZX��ug�<[;�ʴ+�?�Ow�x�O��VaH��u���⽈8 [觙�&F\JO��-�I��TӔ�[���E*�z��C @�	3K�>
�g��;AA�����\/�eԶt���F ���PmO�;�?�e�9A���o�ݣ��'rw�(�bA�֨<���Ű��	T���Tշ�sv"�x�UE��t�=�f\?N���KJ`�2�,5?���9������e)�7���P]�z��S���TAe{���>�{[�NYi��^�;8��D&��!���K���X�p_)����^��U|B��P�8�4��HڄT$��^�)<a]!A�7�QC6�������M�f���t�O	ib<�����?�6U���KѸ�t�k���`�%1+E3�`+1��+�d��xu���}��j���$�L��
lwH��IH�������5�=aݻYH�W� U���;�ꆾ�PE>%�*�hV��"L��L�K�!���3�}�C_��7]P�L�E����D4<+�Q��0�^yX�Un/��e@y͟o�B��V@���k�6�t��c�4�S�_� �!���(V�<��Mhh<s�!�t����$��6�L�¬34��$���!�'P�D��nm�Y�|׎h>��9��ƣ�Q	���5l�^͝˝n����*���M��s�y�Ț�<��JA���zKP"M�Mm���z�7��8�tA),@'S%ѕ��,*f�����^�����Xz�2�P�DT����.7(����e!X��ā����h��&S�����@m��Ra`����G4��	X�����썶p��[��ZQ�0�^G�l�E�����Xi6���Ե��a�"A�t!?���y���C�M��T2�]�6��"z��9�	xA��F��lq �Xx��X��2l�c�Hkƣ����5��3���.�J4��u�Z�����i�����]���e�`�*���A)/�@B;���H��9���9�L+�o�T�����B�f�^~W�I��M2��CZ�L� �U��E���dqM�&4	Ln=W`̮>/[鿜��2uqHQX��=����'�3����#WV���p��Q.���0�c����f�L׆�)ɗ�qv�70-ND����?_���oc�������+�D�5��'����V/��=�ً8��xy�=	ĿY�4S��Iω�ױ[�?��BY7�-�~6��n�lyv�Bc�pȹ�S�W=����t2	����hQ�0�S0�[U$�\���V+����Ի1�`��/�,y�y��,�.}b�ߴ��6e�@����%ˌ\n���,�~��a9ޙ]Ow�!�l1jN'}F6%ڿ�6�M��/��XU����Q��ʸ��\�8r�z݆�?Ӓ��R��k��3R�h>��'�N'�~26P���d�5�t���nL�uj�$g�q����0����E��]LȰjF�X��_dB�����K�w0�Q�(���/�m��y�uQ��V���M��Ѡ`-�1̏��/:��"c1n!K8�I��*�	5U�����l�L��w��x�u�Ug��v���VZQ]\'DgK�]���$�T܏��Zfh��U·�L�E���\����M,-�HӡtǱ��2c3O>�*5}t�SL0��'<s�hB���>H����%ѷ(�H�V�7l}n��XE<����~mx�n!�&��Nc��7����s�b]#_��m`���J�����(�{K�����6p�F����zv�������a������t�l�9�ǍͤUԺB�d��U��G@�s�h�6�����4� y��H��6��Iȓ}��ލMN�95��Qұ,\�]���fY�yA�������zB�I�b&v]k�=5�[�#,�^�(=IjjSd6��:�b�^S�RR����D	�~|��l�* ��!pB��h��9��A�ԗ���E{S��E�Y.lZj�H��-o;�8J� )��gL��$�8���D� ���X��o�?�?�����XL9�����'���Ŷ�S�5i��Ki?�b�ZʑV�Ϣ|�t�4N�<��z�|G�����'ex]&�V��C��#�t���;W1�a��֎�ݝg�/6�[O���}/�_�<
.�1�җ���H)P����i��-��t��Uf���t���.��9t�J������`8)X�i��F�џ����Ki��{�P<��o��@E�' B�H�k�|�?Fp�B�a!���鏟�1ǆ�{O����\�~��K��=E��B�AǑ��]Æ�=u9K��Ǵ�x�3�?y�3(�4�,��B��!H����H�I1�I����r���L��ڙh@��9�	�g�A!:ӱ�]E���"�����)FeTdZ`����d���xR:�\��me2��g�h/���^%�A�Vpu�"o���䉈�][4����X�l��ѕ7��qG�T�zd�$��|4="�wR6K��T.�c���&;�Y��xb��&*����ĸ��1:g>_O��K����?pg������'��:���x	�{���z��Ͻ䃎J,��\Ř�ңp�UL(v���j���7���$;[�/w1/�A3�lQx��������`%�<�/ey��C��_�� ���]r{�!ou���bM�%�Fx+�+��8�K�3�ML��S������h���c��?Ѭ�:�[�7�s�P��Bw�a�I���g������>c籋(tl��W��x�5�^��M����r2�Wm/ @�EU�-1��܂�r�ՐM}�v}9l�iB�P�1_^�ȥ�j�Z��+8�5�kW�5f���!����l�վ�ǃwZwY�eB���GH�%���A�#�<X�s~Os�s�E�Hf�!cL����l_8���
���ƒ.T�p̶����͹��UN�}�gߚy�&���%�F����Ұ^�Q@7̸�����u�X�Y����Ũ�y�T_�(R�TD���)u��t�!���	v�9��HZ\e����c[��>����uq��|(��iO!�R���8%�	[^���C�B&H��H/T��&[�/��Gmk�s��w}�N:�c����� �fIrZ͟�X��S�˫x��Fep��'�� ��r$�#��H���Lt�MI����r�ػ�l	���bl昳\�y�.��s��%��a�젾!�s^/�J�V�ݜoZ'
�;o�{��a�!(�MN��I�;J�u�X*$S��#�/BF-��t���˂��cg̽4�y�d����9F��2[_�N�j����c�ź��' �k�EN+:���v b΃��ƞ��,��C��䧺���bR)����]:��DV�2��<j�3+�}��V�/���.�)NpW�����y��G�|��kևю^���jj����"���!y��h&N�T�A��aL����Д��E�M��k�Q�	�ma���ȷ<Hm7ٛ��Oܨ�R��w`��D�yF��מU��X�2ig,5B���Rۓ:e���3p�װ�y	�TFC�otJ���D(Cu������`��6Ԩ6��w~Ϧ���\W{�IT�|�5$\�֜�x����%�l����3n�9]�B�/�[�au�����G��W28ԝ:P��􀲿��dv=	(Q]ˆ�̥�|;#ЛG�t-hw����"�,��ؗ���Y�!��(�+�Y�O/T��Td�c�����V|M�*^�Z�OcJSNo~i�'>��;T��;�ؿ<BF��j�@��.�1,�������l۫��2��w)k�jٿ����Mg�7VOX�)_R�p�<q*��۽��K�������:v�댍>�%)s{��8R����א�
��R㫕�Ɲ,��.��!��t$yfI��y�)�ϧd����H5� y�/��"pN2�z�jF�D�^,���;�G��#�|Z/��q�Y���U����8"���ЩA_E�Vʄ0I��ʡ��V!����c�h^��������9"�1�NS���Rʤ�Fqُ�� �����b'[T�W�)��ʢ_� Ӏ#)щ<�:G7 '|�����&�T)�G(c��nZ|�����w���g�o��T�6�~X##�3�A"�ԣ����%�W4�/���E4Zwa3*�� �T$I@)}s?��_��h�/y�(HߍOq���6V4����r}`m)v���$�j����f,�z��؟�ǲ�XYm�y�est�oLdq��%����x�˿!�Ϗ�h��E��ͣ�B11�&Fء�i��O�%��]����R3�
	�<T{�k���ȭ)Y���%�l!]�-|W�"p�{�AL,~��_�s�\~4���e����{��m��-#v�!����Y�!��{�(��|��&�� W�U�I�nZ�� ����;�������~#i�Mϵi��bfl�-o�>K?)���$�n+��䅴������X	��L���A���nޙ��Ɓ�i��N�X�mk�X<���+��v�;b���4����S��>�����=0��I��@H?K�D��#,,���T�TSe��m�[e:`HX9��E�<�K�@ĭ⅋O�[�FJF�Yp_!I���E���i}d
���qd ��MSD4c��<	eT\*�
<��qC(�I�6��(�R8Ii<�S���w�|8Hi}
sA�CF�|ü��j����_��ܣ��A,��]�O��*gJ_������b@N�5��1d�e�+���M����1/!��f���O8h�)�G�N�n4Θ��.^�tVԬ��C�p�~�>�b��ewK��mL^��Eﳆ�~̺W7��o��j�?� o�F�q�^Q�P)G�=��X.��<� ^C94�5:)�*g�s ������ Kx�X�e0��XH��!e�j4�߶퀐�����Z�ttt]3JfSi�+���V/?��tq���	[&��.6��:��_��o'��->�3	E����N�e�ϫ�S;O��ܕ�ʰ�K�|5�b���P3��rGB_���W�&���o�r$�\!��]���kF�&&�%�'2`��5j�4���E���à���K/di3-N!�'�i�nRaf�;��/���;p��}�����^SU.�6���:v"�p-p��%�I�x\g��Q���G-�eb.�M�Y�'q,���wj�Nb�9il���W����8�1�G�V��].�_��mSs���h~$��+����BS� ����٣���u��uY����@ $j�N����R� �c�\�ϙA3r�/Bv���(��p�d.~���l�Hd���*�?��l<\���?��:4�k��'�[�t
N�����!k�9�`��Bԋ�E�NZS��Z��
�Q��0ey��]�n�UQC]I��~�Y�:���Z�e+���G�z{��BA���x�%a-�����7�,�-{�����>�Sс����@.OQ���"�ߪ��GL�V��Q.X�6,H�E1:�,��?�]��n̔�R�SP �H%vˆ6��eF^����=��W�m��*{#�I�Xb��>�|ĭ����wa����ED�ȫu[\����*G�Gv%*mkΕ���O��z[9���h���tFHy]U�=#ַ�Zg���mVW2�A��Bر4�)��W�tUH =�:vGySd�d�8*� �bb;��;��]���!�6þN�m�D��U���T>�ƃu�	魖�.H)nF��)_�x6���3�
�ztu��vq�(�΅�Y��^Uf�g���o��L����5�����
�{6Y@0��WKc'�sE{�%�s�������� :d�]���P[ύ��\�R�M��-�Y�2	y�/u���D�Q�hW������_�J���bF{�]���>'\��5`���&9)Z�f:�?a����������5C��D��A`2��&������R+qki���/j	�b-��/R�\1�O��m1:����'\YH�>ݑH���͸x�K%��ȴN���pI�khW�Ib�O��"̺�E�_��kG�k�%�����Ô��b�Cz���1J�:z��3N�h��w�{��N.�̮��>%6���(�k��p�HK����ƜgR��gZ�x�)����(�fy��/������T,���e�Nm�|p�v��9Gz���DW;�T΃.R��	feNp�2��N�Mt��\�"���[�����X�"M���Z�BZD�pe�sm �"}�j]6���|�IJ8�:/��t2�ϝ@Ԁ���6�p��@��G[@x�b��FEO�����lo��ϒ(���ۖ�ޡ��զ�ºoNcޓSS���WW����wȧ���Q�F�����⨲���7�����̽꽗E|�bbyxsH��wZ��J���̐�(�O�ͼ����`��]�en#f'J[.v�l���XZ�4:u{Td�8%����ɪ-�-~������]�dLo���2�D���/�B�����E_c4n}b_�=�����,��mw�!�����D=Tob��kj�-�|�>�>j�c��M�d���^r7��b<K<�$���N�p>��3�|�6#� b՜��yጘ��oj��pu���'�DmP�)�<�|i_V<K� C��M�����-F75��3[AC7�%����L=��p��1~��s.4�۴��2��~�'�Jw�$���S��.��E���W�NJE�1L�=��l�x('j�FD�w2d�����`�]\�9��bAg�*z{.���JA�Y�%v�mk��-�w��J�ۚ4Ka�
��y�7���z��[��R_$�s�T]�.1�{��kKZ���{cq�r<�KC���(�.����A�F�`ơ`Q`�7�A�z�+g����H}Q�G��* t����6�R1��(8�~d��������@�@�$���B��q?��7Ñ+{#}�s��+� ��И/�7���������/8q��=Ƃp��u|�.�i����.���#��Z�f�9�@E>ȗ9Z��;W��	
�&Qx]@��΄���<�]�!��,X+{҃(eS+�l~?�y�1�rGEW݆^�??�@cLLP�0$"ҷ�?nrDML��H��e.�A���W!�%�	k������Oc	�x�B�u6���3��k��f�m~�[��'�9�",�x,�����v�q�.-��g�_�c��~��k�"��g�l�}�a����Nqh�x�g4Й@����v+�p���q2VJ����y�<�~�3��ѫ�pM+w�p�B��_^��Ā)WK����MI��I�>�"��⅛���׵$P�>�4*Bc���nL�̎�t�F3�6*@(��C���� ���䍞�|��7Ѳ�1ZԂ�[�_�B8�I%j��*�&���P?YT\��e�L�u�Ϫ��7+P|"�Y���W�v���zx+]�W)�h[�1��ܕ"�����(=��L%����y�ɀA]�OM8�	%q��b2�i)��
����8R���m�V�@=��z�:b��=�s����@lY�
�TR��<�K�`�����`�h6�]�	|Y��|�0�?�V��!
��$n��n{��P���4�㌐X4��R�o�*}WLT�>[�����ۤ����%5 �21�v7�;Y�k�f��@`�J�9�d�Ǆ.��|x����s�7�Z	J�t=fV��5b�;��(Fn��v�;g�@��0qݤ��Bd��;�M����|�c�O��֑� U�@�\,V�d��������A6�z��Q|�ڪN�(9�f�Im�Nk�j7�X�g��M����B�
��ڠ�"�7b��:��J�AB�{�=���ǉ�ݵq����c�$V/��J�pŇL�琖o���$C��s.
�ۨҩo6@�4����sY�Y�2�笭������.w�)��ꍦ@Jl�ݮT�M���ݣ�n��	b�p����t�nt���>��R���.n�U�� �l7�A��a�`I>Č�˻Cέ�2�n@�o�H
���|��Lk)�8Κ��"��}Mڬٵy�1�~�S7��{���\���w��������,4NM�_qm��^>_�U�Z�Y�X��l��~�d��tL_�iUW��w��U`9F�6�����qݨ�BaG��ғ��d�u�3�C����P�6��J�k j����ȓ�kg�����8,�Rx;� BG�������R���B�hm�nE| /���.��SSSN=$��_�b߹w�
~Y)�M�B�κ��ܨ��?/�O�S�s�oZ��AO���W�^#ܒU��3��:������G�fUQ�M\��,I�������-y���%���?�N-Tnj��7+7�T�7�\�v"d�ʊ
1f��v��uS,f��2�o�.;��͠`0L]2���+3����.�B����L��J>i,�U�����/dKA-�v�����B�I��
�1<�^S~��N��=�/à�#��N����O�\����Ь ��xb�܂�٥xP�{V������I��������SZI�g+n��1϶
kҠ�)q֙�]�p4��-Wf�o}ī!��WEs��֌sLE���L���2A�FD�ٿQ�O45���^�Q�L��i9� \Baޤ8uW��L�s�d��qNUS6�JiTgT�ܓ"sa-XTOˠj�L�@l1�VH��	)�W�ΦD۔�/�lu�U���i��"4���SB2})`y�Hl���Bc^V�<�cpJݩ�`���}� c��c˚��7�S�BI��"NU�G�\�VQ�E+��C��D�e%�qz	�^;[v�3��I�L�C�q�YHf��rQj�`���z?,���T$&�M^{���n����s���E���B�]e]��/��}i��\��[\����*kE���B�mcG>��D\.s�H�����P����u��q�mAܵ���)q����-պ�M�����q���TP�;���ʝ�;~���)1��)�%������3o�֐m��}����#wO�L��� �vT�~���		��? ���l'7�W��2 9f� �4[b�z���)%ԣ�{I)����� �@]��#������!�-���J��c�+�%:�m��f�(ez�ߜc�YвV+>���s�u�fn������I���Ul�P�)�ǋW��賰_�2L)ʵ��Q6�Ax���gw�	/���M���C�ݓz�L�S�'�x\r����×f�9�a �Q������FC"A�N�b{�=��M��`�_*�eD�[J�S��Ԁ�Vdg��9) �EG�C�ފ	w��eAF�a�I��!��� k��35c������D�k8՗	R��;�.��b�ڊ+rrl�Р�
	8?��g����x�@�)Bl�S�N8!�?Lѕ�0C�Ĺ>�KN<����x| �� �+^������g���6�M�Y��0Q�����we�Z�@�0�
�yӛޔ�w���纍���u��s�'�9�~���W�����`�����1xŊ<��L��9�Z�^~�Eu���r��}��Ҽ]O�/���ݕz�V�wݞC����Q�kH�@먭�FO+�� �#������/~q�n��D��Q�
XVҳo�]��Z]�r�E= zjq��1��@N+c�� `F�S�=u���q9��Zt�����O�Ld*uۉs%^�v��d���Tb�Mh�Ü�!q��Q ��m�C��0$Y�\88����~zf�_|q>�{�J����ʤ�Y& C?D&|��_����Ȁ� �q��B��b� k�<Ϣ�Qv: �C����_�>K�<����`�1�'�@�K�ӷD]�<�(�L�����!v�$ �Fθ%R��aׁ0Lx����h��=5�gR�#*=ݩ�ڗ�w[c�*��2r1mrT� ܞ�KePpב�ȱ��S#6#��T�
fZO�0�3U��t�i*���L	�Q*�ؐ�T��
�#3U�3�2��Vj�v�H;Lq��Id7|����wU��{�Ȅ�n�^�|�3�fˆ�@��9�����$�=Lլ�� ��3����͟�ɟd��������h7���p�'?��p L������
�I��rl���r��Z~ٯDCv\�HƫK�2+�`�H��"F�dR4���Mg��9ޕq|���s�,77���'<;�Bݩ��|ڴZ�.�#��~��[7ϫ��ݖ��&s[ޏ�]�)I�49NOdU�21�����kF[��h�TH%`d :�"L�LQ��Y�:���0�9��t<^GpSs�7�8E��c]�n�Yb�f�L�>��U9Ǻ�םj�Z�2�O��3�,��M ��h!.���`��:�b�s��p�3����&�L�Q�����.���Mٜ�s> eyZ�O$��K� E�J6:�@���;R�%��Y�83^)��Z:�xvC������F����\���rD; �9G6ie�����t�v�:0S%�6�{��QV���e���eW�C{b���vU���d:Ʈ.S��og:��:y\��V��} 2��ѣde�X�W�.d��	q;˽L��i��_@f��l<�3��,��9ޫl��g����8������Єa�0�hw6gu���~�j�e��z���-�	�@�=���.�&6�@]M�c��ϻ�p�C��e����jh�:�D��||+�����j�[��s��Ϧ�(�	�o���|*m�
ǲ4�5<���'\�����#9R*3ǃ�d�ѡ�wesmw}q�pDs�����ɮ��+����eH"�>��@x�W�Y�欎�������m7]�J�`ٲ�/?p4��4V�9 ���ifG�*owꠑ��iL+�a<m�	��ɴ��9����R�w�39��X���Fd����9��3�@����+��e�Ɠ�{v�Fv����b-����J���m��I9n,���~�}Fg,W�]����I�^$�)^�N/PD�HA�qz'���1����=��bW�^f��ٛiVciP�-_��h���>���y噒}(Cd��i[ATPҾs�/�jH��r�w�R�Rc9d����}#�R&%>�,6J;��V��?��q��LR��Y����O�]���p�#�n�|�p^���1'Ǉ��3�&G��:T՝V��S�q	�g����f�i�H�S��2�3�g��_�~��h�ZM�:y�v�S>��?���.�I�2�`�{3p�vY�q���t^�R��ؗ���<I��x	 �|Wէl<�|,K`��͑��s���f�`�mF0zw�R�̺u�N?��#o�H}��ʲF�	�� �մ��E��)�^RW���E��hd��v��Y�x�*�����r�:�SnU�~ou�V�G0j����X���#j�婴���-@Ff��;2j���Z�M��yO��+���X�0������3<�(�,ʤ�2�7��U�� (�-�c��s��n�|�p��ㅨ��2>��SfZ��y+�G�h�܋�1LE)BQ>j]�u�V�G���j��"�+�ɛx�`��f�
|Zw�f�<������FS����Rw*l��L���7��T�]�����D@x�:δ���f�QS��E�7c��]��}z���-���c�N�X����""A���N�v`�ʲ�x���׬YsZG��	/������/oo��;;��c��Z��<FR��]5`����`#����>d&��d!w���ޛ�Kz�����=�<d&$@�à>8]8W88!��H!�	(I��4�� �E�0	����9W�<xQ<�	��t����I{���ߪ��~�vU��ݝ&���~�v�7�o�w�����w����C������Nސ�{��4�?���u��Vq2Ĕ�|6i�B@��^����`x�&.;��>y/jy>c|v�t8�s�i�u�F(�Lޙ�Z-�z��R��J�Z�>z9���8.u��aWX��b��vw�*��6\)�B��w4h����� ����;A��ױ�;󌶣��+l?PF��ڽ�a[)+,�x��ږ7��E[�X��$>�P�U��;N���p0�r8�AaP�;��fo�?�~%��ˤG��L��a�e��!�JNpƮ�jc��_q�[�V�;kl��OW4f�&wD�I�v��A��{��M#�+<�Dt����r�2��xm��GOS�WG��6e1�[�v���	n�;��C����QX�������̵��8ײ���SO�N;�����9�t�DHT#��6��T��z����2�;�t�q�{sv7IPt�YZ��M؝��
2�����בN���j�2��x~l_;{���t�lo��{rڹ׋$"��*��vsH�bt���k��*�����Η, ��6]�f��ދ���G�T�h�����L�jc�����O���\����0{̭���?]�i��ARw��lg�n�j��޿�`��X5gn1CЬT��Y�u1�/�h�Le��.��iԢ"�Q>¸K+լJ����^�J+ѐ��k���wΑ��y� [��,��St)�n&�<qW�����ò�Z�m�W���w��q��2��`�إV3�F��|��<��z���w��P�o׎V;�z�Z���c���!��\/���{Q>�8�]��22m)��=��k,�m�Q)��k^[6(��l��`�,��F#񐱎���^�l�2�Qqb>�a���MY�{�s*�r�HHr�V��r�V�]w�UW�jI�����;n�̺R���Ä+�RzԣN�L���l��/N�H�#h��ei�y!8V���e�s��;BEG�!�d�ܨх�]D���&�.2i��\)�1�G�^�@X#��x}^܁,v>�5���#덁�����An�K��ۭ�y!�]/v�R�ee8?��^b;R'�(Ld��@��<Z,�'QI���c��K��!���ǳ �<ܯA OY��m㦗`��b<��B��s�$>�ed���G�х��R/r�~�oJB��ȑ)K�|^��B@z�AY�s��&c7��"P���|�dL�RO���Au�wl;S,�f�v��M���tZ�Z����v�EK�O|�N*m����q���\5=�'-_�2��-K�{�/��ǬLS�>���rG�0��Ep�x*������������.�hV&�����'S�Qʘ�a!4j�S��m�N��`#;���\��+�� l|�7x�r���y8G�F!����������EcLf�r��B d��c,ovfoԜ�VK�@-���mJ�F�tZ�Vj�j���p)M�v�n�<Q��R��g��ZKs�-&�Ʋ��q��Z8�>�ff�a�A�}�iD�����Bo�kE��s��%
Μ���
��[�Bd��3�+�[��a�ڼ�5�=)r�������zQ^��Pzp�n�Ȁ��00�%c�a7q��wq��{S�uAuKH�	q�l��v�Z�^��˖���8���K��u�KW������M˦V�5����^v^Zw���h�S�Ioy�1��L����l��	����IK47��7�^a� �ph��Բ��z��YfJ���Iৡ�%�G`���q�?��@б�.��>sv$��q� &�|@'Sj�H�����{$\���`��9���2�����K=��d�m���s�Lw�;��� ��	˝Tj�ScvO�4gR�4�j�N�R
L�?��� �K�T�J��e��)�jm�9m���|���Ԛ=�;�8;��@؝ǩG���DFL�b#�=�.��Z8�>�od@Sk�ހ�KP���~a�7����=�D� �;!G�9'�+j�(qu�m�p���ƿ��N23�گ�Z|�%���ʖ�CdO#�}�g��.qv;4�&�-�)i���C�R/�P���duR(�,�[R���sL��ˎ�o��S�{V��I�Ӻek��g�����J�l�9�l��
uD�*�
#����/�A��R1��#}�@�zq*�J�0HbM�9ݱ���0�0�s](#�I!H�����8g�w �IƉ:F��4�ܫ40�IM��Y2���:-�b��#��?FFbor7ctb��Ip���:w ѭ��)�k_��\>@��_�j.����G?C���g���x�X{ww��>�y�/��?.�����4���T�{_�vfS���Cw�T�ו��y�;�SO�e+Ҋuǥ�D-�|`w��W����1u=將����B;#O0���P�7o�^ �F]GF��ɹ��ljp�%���A�w !�ƽ��9�k�17d�K��#�a����e�l���	�-����}�k�@�?�����v��v�n:� y�k�naͤ�$g��@���7�Ŀ��/���u�s6Q8��s���ɓz����IEo��@��D��z{^d�⊍K�;�W]s\���t�=w�]۽s�Բ�43=��_{lz�K_�V�_���_�����D`o��N���@T���i���A�L�l�� [#_(�4�����Ї>��R�1cr�4�>�bg�,��Ʀ�0�j�AS��h?��?�wQ?$����<�0eư1@� &�8�@y ;�b||ϳ��]�ʝ1�5��n�������
x�	s`0�3���9i��N>�Բ�bq���-w(�g���Z�6U:�Ԝە��ܞ�voK��L�4S��wC�dT�Bڪ�Ruٚ����R�0��d�g����O~*�y`W�*2�4Y��obx��{k��`C�Y�\u�U���漋/���+z��&��n5m�?ڿǩ�9~W��N�y��6b ���������}�O�ց^!yzق�~*a�8��>�M��A�z����&������ۋ.�(��+��r>G��ӟ�}0��乭�a�T$_`�7���_n�Z�J�z���.wē6}��t�Mo^��g�n��2�RJ��~��t��ek'�?��?�;��Uw7j���ac&>ӹeY���\v� �mDu%�*�
�qC�#{>9":s��rC��h������p�0W\qE�����2'TР.���h����y?L���2���svW�%�<���tf�x���)����n�|��~���;5�~9p.4P��戈Nw���=3�3�} �ukW�jj�NcWz`�m����4Q��r{&����F�of~�rjWji�]MS�O�ם�Z��4ۮ�=Ӎt��@15�-1?�K��s�zPF�3	�ِ�v�=ٰ�}9��/�D�p�����'�5��0a�Jr��y�X����c�3F!p,&�7  �����D�6��3S.�4�ͩ��:����U^�n�����DٰU��5�\��i-���og��>���c�9����{�2�mL���� "ЋqǲpH#������2����\�iӦ��l�r�;�5۷���]_�K���w��?��w�ȳ�j#�QL���]-K��ŀ޳[* ��>8����7\$a��ѝT�<�Q�A��pܓ�`��@�k;� �E�t��(����.L�Q���t[-#�lE�ar��<��S~�2[�Ȅ�;����� � �lي4���W{�9g��kV�j��R}O�ǖ�س#MTfS��Y�n��@�E�Ze"��Ժ����N�ʊT��Ү���k?��y�� <37}X��y�`�.v�� a��QA����:�������b�N�	���{���\_�� ��7lؐI�2����� �eP@���r?���9���F-�S׀0�� I�B���b�S��(G?�����_y��z����#���1�K��u���;���hh��w�<�v��n�Q/������a I��z�D	ڕ#d�����O{��r�Q��S\��q ���(r�$�����1�"x9����սa�L��U]�a�}d�N6Poh�	:. Lgְ���k�M��e���.�4N�c� a��{Lx:��Yg>��{���r=U�3��Zy�-�$=f�e�<�f��ij�Ҳ�'�fuEy���    IDATjt���F�����;YK��Ls���ʏ��Ud�9����l)�0��Z���u��g��Äq�e�Ev���XU\G&s� �er�~�oܸ1�=y  �F��"���[^���~�ٸN�]���ס��s�6H�ֻ�޹�[����/2a۪�^O*�%c�yb���/]�}�KW���(G��Z�利5I&��G��x*]ȇ�� !t�8�{��g&,
tL��^���Jd�g� qɘ����?������KV��԰�);F9"2�x\����p ��f�6�=1^��	+G �c(�x�;�^O/�[��%�޶�0�VN�yu\^��`��3^�"���J��g���Ք��� �J�SOӭZ�\��4�^��Jiz�����S���v���j�?�m��� a�� �@8�罅N'�,�r0a^xA��7Оq��Q�X�r����BL8�����R�0����~{lSc�x���{�gF�H�����C�0���w���c�0��@��@x �B�:����K������ߗ��q!j��FG�h�DG4��R��b����3�<8��m�*��|����W������?��yGe��ʥ����p�x�2]EA�@@��	;"jx���"ƀ1@ga�(����a��Z9B&� g�#�ZV�a��.1&@8�NV�#�h�y�E�1=���rskV�j��R}Oڵ}Kj��@�5�Քʬ��p^�����J��=:5*+�\�H{�&|mᩱZJ�V�m�Lx���G;*���d���+�� ��V,[�`� ��0a����=�����*`L��Ӡ_�=��<[��1��g w�8�#���b	���w�0�G���g/{�U�~����9"t����w�ؖ[ߴn�֗���3��!G81�z��Q�T��dD��3q|<n�F�h;�c-ch	L�0�^A��R�V!��� LF��C�T�`b� ����
�v��d"�	kP��Y��݄	�LN��	+-��9�L��}r��4��)�w@���v=�K	
L�e�Tji�UK����?�µ�go�����/�tA���$���~X�/��E9"�	c�Q���)DQ��Z�N���	s���Q�9By��F�҄#����
��Ș`c>��h��-�&x�2?䜋a��r&}����Z�HȜq>K�;D���> �D�r�R�0P\)W>�q��Y2&�o�r��mY>��	+G�	�<����y�Atw�Q�o*
ed�a�0a�)uc~G��	#�S��-��&���l�P1hX/S;��&L��LX��r� ,�	�	�|E�ӯ�<� l]'�# ��R� ̵��N�9p�/f����l��gow��61��# �j���s��m����&<�A�&	O���=}�SKӭj�:�4��ѩQ]���X�=3�>�'�H�wޗ&�*Y
�kD�]�y8�� ��'抚0Lx!�s�	S�h�21�u��"fg����BrD$&��RL̙��? �L ���!!�� �=�	�Y&�g ��N���	D ۧ�=��Ȅa�BB��	wCtK)]�eo���x�8�kA
�_6]��v獗��~��k:��r�!j�	3� �0#��ZL� &���}o>o� ��R����f�a�R�Q�U2�Sa$�\ef��n4A���@g6�� �L�Ɖ��QR�����K�;1�=r�W���R��+>w��$%���e���_si_�/�gz&�zr�Yg�t�Ks�i�@��4^n�rk�|��	ۃ7Y� J�SK��JZ���4���ԮN�F��=����O\�vݿ3M�Є�~�8���]>+�	AXa��1���A�w���0�	h�Z�����W�l����8A/�&l�@(�/@� P�/�cC}�����%��`BX�K ��=��RF��sW�ƍxi��s�� a	~���.��%�n�d��7�}�D��Fs.k�G�X�k����w�9/֨כ$���>��E�;l���S:-yT8�'0�όV�D�<u����9Y�a@
��B Lc����]Ӹ����;\��o�9���c�+j�>����\ <#*�3�%��;�񎮜#t,+��,̆�}��O��O������"7�w�m}h��c��@0~<
���Q��� ��^���k�涛k�s�=���H�֯J�V+��{S��>�:�T���$=dI놪�"�Zf��jj��Ӳ��R�6����|`W�����������R�3.�E���6�J4�Ձ�� �ع瞛m���f}��`�=�~�d9̫@����*^��+%$J}q��r��r��/��x��!MG��^q�_��aꎸ}"���g��7�pU&�|@�Uϕlp���:+�5}vA}��_�܉I�&�ўMF_a�"��[��Vf�JLeT�奍��L��/a�s�  ��+קs�9{�����F��P4����T��K�g*�����6�����??�Ӏ�Z��!`иѭx�k�PG�<*�5T�����p���x��v��m�c��ѹ��+���3�����q�����3p�7#��z�wup�� v:	uI�v"�r�,�@�R�B6F@0�7��l厲wzw*wHu�L%�O�	JC���vzrn;uJ�t��.�)͗�?$�I�����gg�\�,'�!qζF����开ðW%7�L��Ja�Gam���{�mhk��[��`�\��z\�T�s�|��U��|����+Qh��Sڟsjȁs<��(a�+'�B���;/ u����_�k�\�?$��B&���	��sR2aޕ4)'�f����	� ����m��ǰ�{�	�G߻�es{s�	�	Q�'W��swo�'��< F�ȃ�E�Ӈ���z��X5B>�|�+�7C���Dy�T@9�YN�`�#�tw E����BY�{;���n���\~^4�c��5*#8�g��c�%ǚ��e�<��kG�<���,Nf������ێ欲J��;���r$L5�X�2Bml,��͜f2wn7G�3(3���R�CFo��vE�[#3[9uJݝ���rg�Tx^K��l6�� ����9��;_!�[��ڹgjF}�,g؏	��I�eb(	H��r�e���1#Iq�s햿%�c��R
�k�>��@�}�Q��s,�IP���2ǵMٵ�9��dE�"y�
���s� �sAl�ޭ�'l�믧�a���.�b�'\��u�-7_�n��,�OS��e*9���5��;�� L��
$8ډ�ج�4L-�M������H�{�~��,��Ÿ�[2p�<�09�k��w��ϡF仃�#�����������Ռ�P4b�se@�!2x�`Y)�@�=ޭ;����*j}�2c�Q����dڳg:w�����]�_��J�(l�����xNi鋏� 2���r7��lf<�̴�e��i�T��;k�ژ:q�|�w޵m����i[��AS�4�^+�B��-pm�%@�o%��mS����$]}'�<���8a>,�K�����9DGy c0c�/����"������[W^.��PO��sb��˲�񪫮���SNY���·�t��w���>}4 ܨ�Ҫ��U�ze�#����Dt ����o�v�cX�#G@�u�u�96f���e��m�y���hn��Q@ΑLY��y���)�=���4���"��Y3�]�0��s�G��2;hɠbB"�*0+KP&Yב	��b�֭�
p��1��m�x�,GĐ�ٺl�,h������>l�=�z�}25�����fNٓY��a�|􈔥�;�M�eE�q��H$M=M�\���i/�BU��{��s�;��2_�U�e��-Cq@�?���j>�y�s�9'�>Z,Rk� n����\�} ��O��&L}�f����,��d���F�	��c{u��+����3�8c�bLr������fn6�9N��/H��N���{`>D�Q0����o�[��u���+�뢱2�����?�gBۘ���'?9?)%��9%��&	���$`iL\�g�E���02Y��׭�ÌP�Qɂ��80(?Ȗ�`�r>��f"�y�^2�AL*{�;�ZwϹf���c��ɚ-�h���p� A&��[���;ώϦ�e,ԩw�F3U�D�/�AD�0�M5��Ko� -KS?��M��ڢ����� !����%l��%)1.��t۲ľ�v'�U��k��/���,- E�s=�(̗�)&�ɦ��+�����,�L�9��6�tؗ$�(��L�{�b�6�1�ܰa����~�]��<�>��n��<@xl�����E9�<�����֣̄͢��i�bG��#3f�W��ys`\(��a� /�1Ǣ;�-S�0a C��VrԈ���s-�@wD�����Fg��*���!���6��;��\��VR(x���a��L����>+�*���@�� �����x^|��k���|4��֟ݎ��N��8���gV��:�%2�l���}麉���C�8�AX�l��HF���CQB�]e�\_�I[��;��l#�g4�'��{�����ne�[��]I\��,_L�ﵰ}u�P�c| &���|en��}�c h��|�#�޽��� w�'�-��IY�񊃟�籜��Ah�!��,j`���6m�t�i��v�};��B˄�m�㼩ٽG��*�	31��lot���y�幹�A�҅���ő#dt�?��2aN cbε߄��b�fA��1�&�*�@�gu�ڭap2z��	|�}d��!:�g�3�\�<JCq-�����!"���xΑ�����!$�l�=J9�݂z�ϝ'�z�1 �;�ZBjH=�!�,���Y~�)�~�VsS�a�u�N��+��h��}ɬd�F���H��.��&���Q��DgP��^Ji��z�����w�C��r`'j���g��{>��ًz���JH�>��d��k0Q�¨�<�9��!I�I��)r�zDB �Ω���[Ǒ�Y/Vγ�l��ԽK z}������Y�����^��_OG=j]�7�R9O�,�D��+��y����	��0q'��s����x�.�O�8�1�]�����OF�ae��N����j]�!�ݒ����Ч���9�#��=�%�3�D�����' J�	|�A��'+f���$	��`@l19�9�9���A�_mI,9��7H�׿���9�����7.=fb9��LL�q�?�*S���Lx��`�x�1b��{dc���Y9�	��^3�?�����+0tm�;�Ły�\��
��`���l�N����?�:���8�4��Xc"��D��`�C��8̤��_�vԉq�s>E�2HT��IO.��M�6]��r��w�ly}�(V5�	���W��g�˫�ƪ�AX�(6Ha'�tK��t�8b�����o��[���ԣ���[����} �V"�l�8���t������9�> ��~�<�w8���m8������E���?��qz�1p�	J�?"&8�����b=쨕+'z�b���w5��u���Qwo{٪��Q$[�	��hPմs��4>9�(&ܯAc��j�`�:	e$��ް�aF+yn���5�����}�0.����}�5Qx�R���y��r�����#��?N��	n�6�M��~���\'���W�XLTw1�I�-�V�W*���#�m7�q��-/[��G��g"��j���6wg>��n�[���̣>�䟫���1��� Ց|�{�a�H��s��j����`<�����|�����]]w�u�j`��������Z���A��z� ,�ᤠ��N"F�̶U���,q����	L~�zr�W6n���%�# ᱻn|��{�z9 L�V�� a��L{oγ2,Ns�0o���9���+��V�P7f�~?21w ��=7�n��*�v�;��v�wys���q�r������a��;�j�+#�\�m$��(��|̓B�x������L���x���	��[��֗?�)O!��ȯ��,���nٚN�hw��Y.�(�u3`��[�,�s<�ai>Le�����1C�z��O�3�ar�~����(�@W&�pO���y�AL���_Gd�Ca(��X������g���ԐP%�w����3���?��������֋9�@��SO�:�^��A���ׯ�~��W6�fb�ݖ����Sg��[�D'�%,6�ofTn�+��=��w���T������[̳<���P��@\�{~̝�x���=����l���{��#g>���R�[c��,=Vف>�*��t{@9���k�S�ʠ�)�r��7o���SN9��Ŵ�� l��r�ZjV��)�R݅X��������X���`�����KZMFjK(���[��:���P9b1��	ˈ��b�q��A���\l{ŕ'��+5e���D�$�i�{e��_tԁ�ㇳ5��`��A�\��W]u�yK�y�ܭ7�~��0��c� �q9ڒ��\��s�6� P+��$��A&2�f�{8�ȽnE � �� .�D�E���8Y�jN@��f��u�����)��7z�#	��M�9��;�a�Z���j�Ì��uy��/���F{;��v�#W?R�k@Y��t��#K!y�@Ў��
eCsK�7y]ȯ�>+�Ҍ�in�w��E�nQ4*W� �,q$c���0&���,.۞�(��>�F;r�!�m\F���6B�g$i(Iؗ`����0�o������谍>�p��(���9���(�H]=L��+f�1<�p�d(��G�ɑXd�Er/��! ,�XH��VJF&`��y!σL8I ~�0s�-Yt�#Ev��8�r��0� L���y����g�0,@�\d8r��8�5Pd��0L��~��v�1�v�>$�1��c�̎7l��VaE���U#$GT*��]y�/;�.VZ�ճř�@�`�	;��	�9+G�	��Ȥ���!�mGnv��� v��y�a�h����!Z�u�
�醝.�$� \.��f���K'��	o}q�?���F.�/c �����_�żݒ��ѥ��@8.m�G@xXm��P�@�s���� �0a��[��;�dA�/���~�����!?��s!D��k��D$���	Ah��u2�c�ڞ-�ɺ��6&H���5��r-�0'�L>�;������ƖE�^
͌k��刻����hd�<�Y����[���y7�
[���.�L`�bbr:>�Ƚ�ޛ�u��s}��VH���7�t��`�����{mٲ%��|��e[,⹑����q9�^�B�R�~u�,Wsq^\��O/-ڰ+DM@C�L�+������ص[w�)�p�B�MxII{p��?�Wd��X��.}��gQ�I�e۴;OOH�LܐN�ܾ0lb����b�PW�@������'��S��T�KʱI�a�&'|����`"2CGgwדN:)�b�c���W i\�]��b�<��>��d�@��k�f��ʕu�����Ή���!7�i�������H?��?���_�%�n�S����1���V7vV�Ϡ�f����|�K_ʠ��I��^���];{�3��@�\}��Y]�'��C0����֑�� ����]��^�i�������`��D�;�=Ԍ�e�
<ĸ�2[���g�gyt�W~�~!GY�C4��5�{�����ڇ�T1H.��}�W.]�G�!��H؋���җ�4���+ۨX�	&�C�@0�������{���
�H^�WdVH0�w��]9��k���N.����Q��,u�cZ'q���԰��ߣ���i�π�Fa���.|Da�,z�=��[-]t�E�q�{\�A��g?���c����3��_�u����s];����w `�^�'���9>�{P=Yp��r�D�@�h���҃���U����3�*��    IDAT�SG�`��8�/x���J��|����y�>s�"~�gӞ�lL)�q�^{mցy.�����y��;+��>�����g�4�m��詍b��# ��L��Hq?1ȗ��e�	c��: )c �aN��3t�p�]�I'g��a\�}�{_ޠ�� ���
p�U���5_d'�Q��X�����2b:��Yf�Y뉎{��f��D�'�k�젋����~^��^l�~��s��l����[7$m
�������K��F�SIF��͠�WN�j� 4H
�*���U�
S��?�4ݿ��X����yW���-�{CD(�r �F��`�\�m�b���p ����R~Ҧ��Mw~�����������?l�#��&�@���8&�KÌ�&Ʀ~��adweS��i��?~�{ߛ�p��T+���<kT�AF�q��s���b���xc��S�_�T����Ox�2����:0&�*r Mg��;���5�I�y�c���|�A�B�zի2���������|%��;U3�������������ۜ�Q���m��sd�QۥLN��[���ҫp�,z9���l��MR�h������1�K�,~.GVjRb�l����� �̄'óAF�j$:T�;<�6X�s���W����W,Y*�G
cl�L춊����g�O̩
*���B.Ԑ�_�,2C#G������<�Ą@� c9�X��ʢ� LP�e��b�D���c���]6���>��Ol�
{O�e�����ԑ�鬀��/ǲ�9r������=���;rė���<ؙ��zg��nY��A��p�a�T�:�5~�9��b���.�E;�����W�-j�Q��3��('0/������� ����dFy��(q��w�v������o���F���Q����Q䚥�Q�5�K��W6o�|��S���!a 0�3�8#��I��[tCuU�����	�2h'D���p���ja\SƸ�b���9�=a�L���fi��놌�  �����0B��VO�s:$�#�L��(��ZL�!Gp�TF��L��q����7�1�9��������	�V��9ka�D��AH��`xb.���Aח�r6C�Q.��N�ˉ��ROFQl�Y�zV���v��6�F`�w$5'���<��z��ȤeД��2�G��2 ��W��%H���C���ny� &ܚ>*�SN���m���߶|_J��S���f�y�]u{����-:�����Ё1:.���ݗJ4��A� �@t��&�@e!@LGD{�����g�� a;���� ��_��E����#��֕n/�&���d�H	</� +tL)�����6˶�4�7�	�3�r���|�#�,_9F@�ikt�8�[���A�?���@�!��O��Osx���0&l=�~�!� ���w�3�atݵ�"ip��	�c�a< �w���k�ʹi��	��|>%�v!��y�(g|^�A�;v�P�n�t���Q��K���)���5�[~��uw�q����zXkֺ�����[��jz`)8����{;D�7�4���"�(�p7vh(�ݩ�;uA�c������9��>��W�V�	W4N h�����8"G�(���^���năB'�0l�PX�F�1�Q�_����!3e���o�g��2�
�<Ϫ���������8_�w�I��z-��;� ~��^7�o�+�№�ɵ,'�����p���?�=�FZ���N&qO��>\��MozӼ�<�~����0��'�����alOm�:����7d eҒ��|��w�ˋr	�9O���-]�G9�6R�,��^�[�@x�h��)�w&��pq0u��aus ���#��q��N?���s��<���5�0���� c�} ���+��vw�u��.�r�}[�w��9ǿ)|�����mGJ�ꕢ;�q�c-�Xi�� �����=��j[��O�
>$�����'Ot�aA�^zi>%^/>���x'a��a�D�7M�h�S_�E���l�)��wd�B�:���Y��:���y�[ޒc�9��,�S��L�B�����s$e������M���>��g�3E�0���z�	##`oN�E��{���afۺ�і� � l���7�Xwڅ �'��ڶ�@�����r�K6l��p�{��VP3���/@ ���Z� 
������eR^�cʽk�����0ꅻ��2acL
E��,�����)<��Q"S64M0��ו���F�TQ��������i�2>�z��B��MXu�yv4o@�mܓ�Q�P�����������/Lqnd�z%��Y���M������e�.��V�ݍ��H����as���� ?���̓�� C癉� zV����� �/|���$��~�_�'e��X�\��e�FNP��x�esPs.���Z{� �ddL�2X�p�R���.��g�qƶQ�b~pZ���7�{��;o�d�џ	G~�]u7��~S��v�0 �<ủu�
���S���;��;~�Cc 0����ig�`�w�V.g�3��Cc��I��θ�u	5Z�(�sm�=d�~��p�m�96���&<��3&���=�L�byY��=#X<qp����g?;����E&\�rw]ڊI?�vA\p�-b��vRʲ�@�2�6���^a�0er���9F�	����G>2ow��R^�-�ﬣX>b�#s�1�q��5»�6M��Q(�EmZ��kDy",�	�t� &���/��U����2[���Z��=����v76���Zٓ%`������J�c�k�ޣȾ�u�N9B}K@�5��0&�M&�p��H�x�f@6�������91��5�(7X�β���Ŏ;��
 Qޠ��� *���Y��9X������ d���� ��>�R��(j�N��J �����tz·5��Q���D��v2l�&����4��=�}r<���BR�;��@
�E[�ي \�+m�6d�!��'a���g2Yf�*F%$�E�*���]>A�ϯ��W�r�)�c3:�y�5�&o���AL��Z��
�$� ܝ�|�+�<R�I�n���N�Eᢻ!$���H:s���81' cp.���u�00\%��_��_�bp�Ӊ0NB{X�E�b[dg�9�Y�As�E����ɒ�D����Ʊ#PF�Mt������B������H g�yf�>�Iy�s�o� A>@X W"Xhb.��I�a�`;�vއ�b�+�㱄�!GD-1u��X�GT���g�-���@m�m�M� �d��0�'�m%4A��9ʤm���o��v�hH�� ��D�8����H���t��������HbJ������]�� |��/Y�c��與��0�l�{��[W.�N���I\;�n�t�ob�{nT�=N���ӊѐ�y_�E?�\Ɋs��jT�\�E1��b���#�.X�����ר{~��pbN�j��a�]��D�b���=��
��6�hA8ztN&�.����y���vz�Z�' #�������b]3P,�JF�MqON@��cT��n��X�e `b��퇁���֊ \�,�w�S����@��)}d697`���zaĸ����q1n��1@�xk0�f�&e�]B]����!%�9Qk���H�r���͛7_tꩧ�X��f a�3k�����ﾜ���D����{g_�Cݳ�a��h���}:�����j��0&�TV'��*q�Y+�K��K�cdE=�:���lK0�1.������jpAR�s��Nx�%�<(b�덢SzO���
/�0,�C��xQ�Pg��4`���d)��k��_	��Y��z�����;@�v
+���+%Y*�Y14[!��� ��N��z(��я~t�	��j���I�0:�y�hJJq��0�@38Q��-���9�F;pMV$���DB[uP���,�%�L��Gς�2QI&�G�&������}ǅ+�{�2������y��4��[*wR�\�����I�V'�:�<�Vnw�q�$/�
��o&�*�@�\�{��{3{zI�&�D��d�2���'�.ty&���ҁY�u�)�dŽeb1!T���E�w�f�����	1x�i�e�:7�M��1�î��w�Ȳ�w��璙��YR�ַ�53,~0p��0a��v�#�EpU�pr���dH䃞�`�nɵ-�sB����wK��e�,�!Ә��� �P����l��	�"���a�{���/�\�R`�N@�� �0���^i��IV�Q�ʈ��<�fFك�x,��wu�hoJ�@XFo"F3��\2�'�]�s%�+����磤R��H�zR |��͛/>� ,3E�貔V�}�4��\�䀵
����I�v)e�&�H�q����ie���S���Z����P��*ai�(�`? D�Ȅ� l�f9)#?��w�x#t���5��X���k6(uS!g��$�J���X���~@c2t�g@��{B�`5�ıL�8b�j�Q��<h��6m���O���~��3�p�,���gC�ޑ{��@�7,�{�"Pdi�8�� ��g���F����8�F#����q�!�D�VV�#��aA��A�:�^��#|�E��BC�U6
%�%�� j=b�Lގ�fc��v�-��ǹ�؆��͹A7����=~	G��:� |���ޣ҄�j�0�vW�7�r%�sY95a�N�u��*��\��.�J�J	�픺l���J�fbq��u=v���iPf�k�u��s�9#t}�������P�<��2��������s�=FP�ɢ�s d�5���\���ʬ�	�� �`����������5�&y�8�Ir<	'�;N��=����H;7:��td<��;qT��Ǆ����e��´1e�A�|G2(��y�����[z�ߜ'���Ǆa�k�x�`D�(��ނ^	�h�
!��KY��r�D�$G�������A4z�=Iw��2^c�9`�|ꌗsD�� ��R�t�[��֋O;���E�}A����[9�m˥��c ��Ċf .������ۨTS�\jͤ��z���U�ͥ���j��R�6ݪ��ک�.��c�fsY��^S�7V�z}��j-�t�Sc)��J�TM�TB�贲�� > &L�ct���/كF?�yR�mW1a ��LP��bd�fň`j$����0��)���f�ê�P�� �b�ѠF?� <��t�g�m�E���a����ׅ��ѝ�Y�����,��5�r{?����[zP���_?�L���y'�9�Aa���rϵy������d�9�LX��!���_�F?��p�~؛Ǒ!�&���'�<ϼ�&H��p�$h3�.H9鷐&���N�T�ߍz�9��c�)��ฟvUl�C��o�d��;фd�M�z3W�X*�����J�Ԭ�{R�wn|�����MscS7�'&��T���6Y�ٮ�ʹS�\i�&J�63	�+�����ޣ�ssO*��=��nWm��U���j��J\�ԕ'F�$��\Q���?��Og��I�/��8AӑV���NZE:SV���w��Y �(p��>�:�VC�]B�Ыђ18����Q:���֋L�2z�/���(.�1M�ɐ"���m�l{�e�꿾`�C�*G ���w�Ű��ʄ�7��A��0<@�d&LPCꢎ����Ya�c�鉆pBU ���٣��,�~ �@v@�brv�&̱ڇz���ԍ���^��� ��7e�c`�����AYf=���r�|ݦM�^��L��0��#R/��*����oj��Vj����3c�2�l�w[+W�C{j��Y>v��욙�������l���}�n��YY�L?��灧����(��i���q����J�N3�6�r��A�A �+�8�!Q���vt��F�㊑ZQ�R��+NRq:h42��������t��R>@�c�"tQ��%�<;�2�RM���#��Rl]�y츑!Z����o����έ{�K�ee~�{�s�m��@AX��>�iX��,�\x> ��:wlìuF�D&��h�L&DT�$S/z%�����`)��S3p��})�3� 9"�Dz�1W2�0�)e��[.p�D�µ�b��X�QZ�m|؁pK+u2�e�-�j�����Z}nrrkk���[��k�+�];��� C���sL{����v�|Nm��?9>��G&���ƚ�R�MN��#h�0#�E������w &��$KQ��;V�
V���t�4ѫe5�R��</�	a'k�+�RcVC�%)�𷱿$>gԃcdIԝ�9v��,���<����@A�瓝Y/� �?�`��	�3�fT���E&,k\���sBNonX�h�1�@�a����)<��A �|��^{2���h6���Ɣj"Qq��;X9��0�&��M&�aÆ�O?��{c/5��a]W�8Ƌ>8�e3��TN��DjW&��Junz�����U_k�\���cn��导c1�*{��k�֤��k;����};�;���g-k6�[֛�sqGδ������R'�zr�Y�Z��7y�n�����1���*�#'��D���iH-����$,� �� �l�D�;����Aȴq�H���Ag�I6�:`��"���@eaN�EmW�Q[t'רC:��2�������v�(�Y���eT{>P��� L����'?9�6��N�pϨa� ��aϩg!;�͌���0�{�8^ ؊9����Fn�G����w�oQ��;�x�T����<��?�	�Q[R~�;�xE���eMxes����!�{��H�r+5R3U:ci��2ͦ�{VL�6�f�[��]��1kn��4�5䨿�D�����{w\���Ϙ��[1^n�N��J�VjW:�A^��,���8��	'��9�4^��R����j"|�۷��]�y>�0��D��J���غ�46Q0�h���,�`���t,�����Дy�A��=�fmٸ�Z,���ۿ=����]��g"K^�u�c��.�o�狃���<��|�8���\�B�a'ƬdQ�����`W䦀չ��kz��e<�4 L�.��zأm�u�V�G\5�g=��*:��qo~繹 <L�o8X���L�)C���}j1vd��k&t�&��67�sD��y��{D���.���Oz7�����p���So�;kd�4�\��j��i��>�N�vܳ~�����zm�?��/ݷ�وv�c/{׉+v=�S�������?eyj./��R�B��f.�xg"��Ĺ��t��Ǥ��>+���X.�fi,����H��ܔ+C�m�p ��  �Ah&=hPFm&���=o GM���T��I8��2�  ��"WL��F6�� t�I����l���΋�శ}8~�7x�g�,����3~����j.֐-F���ڪ� `eY7;�,� 4�5�19�Xr�m�\k!���>��e��c��q/z<�����(�T@�6����C���84D��I�e�<���LDr�����3�YP��>t��҄#I`��J�r�[���2nV�	�ҷKS��9�5=��o�?z��\��l�����4��������{�}I��/XU�?�֜��߲�I��zf�0��]&�0��t�G>�'$��Ս�8S<�9�L_7FL�.�/��Ĝ�ј�)���?��?�,���.ai�u��0�0����1�W����y�%�X�Łf1 ���C���!Vv�le>G����$.3e�! ,� 
�w�w�k��q�@X ��q�#�u���X^m,�v;�G�_�d� h��I{��/}i�&��	pрIlO�RJ�@�X&'m��<��B��2�,޹���t:��箾���<�IOZ�dµ[���vl}���C�0 �3�U�i�9���c���=�c;O\����E����Sˡ    IDATuO���g�����w���ܞ�k�Vfó��J-䈉�x�� �1I���K�v�ַ��uV;L�C��#s�7�1\:�
�$�"�������&��w�+殺�̘.���1�����}�p�ا��� v"ʮ����-/E���^*-ulb�&7Dͽ8��"G�Ar,2.�9)�"��f��d &�ꫯ��a�N8�	�_��_���ш����)��@��E�������ZFuv�.e/ًԦH��	�n�5��3�]2�'M��wd�`�Oo��Qn=������yQ��7(?��uѫ�F�\���͛_��'?y�bl�@\�L�����̊�U?�����w\���`�}Ҧ.�=p�oMn�����=O��'+�v֨����X*�K���Ǆ3�k¬�۽����.ơE�"�L��;'2��8�AV����a59�.$@�}��&���4��t�a,8@�$�u��`i� 1LV�N�*;n�$�����8�?G�T�81����O|"���Q��y��8]H@N&� s�pm[$��l��F�j!9�p#R<&b�4��T\%���s6��jχ'lzMm�� �a˖�3\���Nˀ�4!�'�F���d��U������?�R���96�E�V�}vÆ�}�S�z�blv�&|�^�~���1�Fy.'`o��Sg�q[��{�Gw�]s���z�m�)����+�����tѲ���c͙��R'5K�y&�E��?=99rX01���5BfE	�2{�����(�N�ڀ8��!�Æ��"󛱔�� 7 Lg�%"���Bg��$t@����7��ܗe� :PM�_��A�p�a�׏�.F������u5�{���|�DD `$��%�6_a+L�E��k-���Uc�vŤ��7֕2	�c[\C@D��w�7`��`�b��=J@�rp<�g>����lX��; �@F��,V�Nd�>�&#k
v�R���ƍ_w0@����c�s�p�6-k�֝��{�9q��z���nԇ_����ZsԶ��M�}׹��{l<�K�k����m��]��DG�Kt�**y�vޝ��|��&�F,S�9Y���@c������ʯ�J�<�){n?�:2\-:.�K�q��=0a�4sNx�X��v���\��\�t'6��	�vu9�b��R��b���������mʅ��>`	p�l�� `NbE��u�Ġa�F^l<&l���@*d5Rx��a#8�	'�'�&�]�;֏�� ��&�0���MS%�]=�kRâ#�?�  a����Rٖ��x>=Fۓ��n)R�0O�� ���/��u��~����Q��<uPm�+��Єg˕�_w����?;}�	��c�E���n1�{�M�NW�?�����w��̩V}Y�4����I���p��/��3���cn�@;;�Fvg09����d"֗s\ygG� l���ς�7,�侔A���PF:2�� V��z���5!G o8��/�����l����\������&lG��]����8]��O����*1ۈv��`��9`'��� ���Rmu���(��?+:�Sb$�ep���\ĳ�l�76�A�9S 4���3�F��`�7eP�Xj�� LY�YڌVN{��K6��L� ��\�n���l�0 ����]�nH����������2&x�
~�����۷^\�v�]�G�*�6S��]B]��4ӣN~T:��3�X���������ǚ�UG$؁U`$]ѭd('��e�'ٶ�`�%F���L��c�9	;����G�e�^G��xc7���J�e�Pf��06�}(�0H��8���a5�خ�\�Q�})�sr�:������N��8qE�Xǃ���; �$��cӡ�Wd
0�:� ��[̑A,9�n�),�KԌ��
���@Oe�����2p��;@��q��s�OAI��I�H�-A]����b�Z�qP�+��"gt��w��kq t,u��9�6p^E�W�s�R�37n|��1�Em���,�0�]�Zz`�q�O���n���_��Qz��9eӻ3q����ݵ�7�7gO�V�v��*�+�Jn�N:!��ſ��kci|l,5���j]]�����t؅Ҁ�vtB�	��N��g=+O�D�Mfg��}��N':�M]�T����ݡ�/���� 	�����$���;`QtD���#�-Ĳ�E���ܶ�2�DPv T�z?�C���	{ �� Y�20��F���E�=�A���u�Yy~ ;�z���xGdA�{l���2O��J̮I�)�ڪ��种aĬ�ע���I�r��B���Dw�(��+��Ю%/��mذ!/��_�lk��#y5�����O�9�x~�՚+�˟ްa�	�2L���X{��G�~n����o�C/�1������;Ϛ����V4�>�Rn�Z�.�M*�N'<��.��rs�T���z��#� ]���^0�=s�J��b3�Z��h)c��#G��e�E0.���_��.�!��+�`5,��ED��H�9l���ʈu�`HLb�"u��bp�]�]��n���^d\��@�+S�z!����ds�>�%�� f�2<!@�A�$P֫�>mړ6 �hK ���Cޠ]yw�Rcܱ=mM�<���x��F}p.�b����N,bC������g	��\��B
EG80�\�_~�<�>T2���y�	K�[�"��������=�3��=v�-��z�Rt��^�ɿ���[~k��[^����G�*�Z�=�J���d��M��	?rb:󬗤j��*$���f��r���KC���e��x���
`�A0J�2�	�+�As�	{� ���ɒ��눎�B�saU�J�ɽ`($����` �a��2E�Ƚ�Xb�/A��8�q�g�}��f�e8�m�Cu|�m H�h�<�̗�$܊�>�'[Vo'��m@���H7���w���Æ�x9�c[��@�bsM��͔���[@S2��|HD�@d��v�_<��7�$F9����IN��v��="�a�0w���;8�=�u.x+ō'��6dY%6�;�$�	\�1?�i��A�l�����+����@��91��y�c>=��Qn~��YhZ��'m�n����dٖ[/[37}R�2Smw�R���*>�7�H'������Zᩉ��nv'��v{>�A����LBi �u�d�z����,�
�-��he��	�z)�b�iuDϧ̰6�Z����T��6��(L�g��`��ι��cȖ�*?;�3�I��I��2���D�������$D� ~�^�=Wtw�`�\�kB,���"�]��U� );k ¬zd�מ�� °W��6x&�Źh�xI��sh�N'��=�kڦ*�I6԰9VJπ��EM�kEF���xuf�}��x�����xhw�8�����ڰa��L����}B��{����ǟt��xMw�C�z�5�Ԧo�q֪-��Κ�=?2V�)Ä�U�J*��S���ؓ�����Y�@�hu��;�C`��>2R*�	;Y�F+@�M\�'� G���9�s�F�� ���r��������\�9@�8Sadh��f�j{ ;��E|%�q}&��0�v�������E�+ھ��n`<�yœ�~aꌥ耰��;yw�F�$t��/�b �=�7���t�#���jK@��L�~͹N��,�/�2^刮u���|~���}D	�ߌv��&.�G�C�6�]{��0����b���mګ�Vh��W��a�]��kN�������M������~����7^ݲ����l�t���*ө1¥4Y���N>!�uΙ�����R��������D�B�U��#��QtⅲEw����7���_W>>׏�8~.��,�w9�spY��5�% LP?���� "�ᚬ,lqy�g&FW�]3"��@,��Eh�H*`����3��������, ��F$�����6n�-Ѿ�%>Äq�ѓiC�Y��xC�O.�0LM�g6O�A����,���n=em���>���q��'��O��T�2�~:L�L�v*��se����(Ca��1�uw�y����1�R3�aQkV�s����kl��c����~�c7������<���󸍟Z9���WOn���k�{���S�5��6Wf��&'��U�צg��ϤR��N:�Ĵlr*���lwC��H\��]��6�52B�#)�����t�x|�C�]+v��Y��;:'1���V�	���9�������6��� 9�DB����;�%>�%�ΚG�x8�0ug�u��8�s���۫V��N�2t�Q�G �� L�	_�"�ri�G�6�d�6�@�k��6��b�y��QF3�2������a���Mm�gs���c]x��z��uE�NC������hO��>�ܴS`��!����3����}n~��z	����ʭ7\�~��W�g�n���I����\J�j����c�g��������L%v};���n|��m[ߘ��e�S�z*7fR���J�R����������/����Dj�Y���E�*�a��
��#D�#��{a�t
2_ѱ�p�C/�r�O�C+Pv▉��;�0 Ё	Q�3"W�v��vG}��g�	����/oT�ڟ�^�sd[2E�ⲛ �v�	�c�|T�Q2�����I `r��	S ��O7��m3@��e���@ȵ����=��1��,,bGp�+��8pM�E��j�� '�%(�;.tr��fH@,>��y�������D!�C�0�h�K����
��6�'3E�"`�\�Z���_�t!jh�v\��	��@��Z�j�S�J�LuC��?:}Բ����,j��RT�3����*w�������dgv�T�����Tnv�7�6t���T�=�ݗ&''�o�Ư�����nTD���F�F��AX�(~�;'P����P���x̀����
H=D���Pnf�)�g���Â���0/_��R�C&���D��sd& <�	kqp;��;��j���y3���] 󐛁�u��~ G/	ǐw���c�##�g,�׊R��b�ݐ[�I��3���(_p'yv�KYB�r�w�Q;v~������}�h�E�1��z���Qtnq�2��ā��Bl���~Ll�T�@c�Z�N��Ax�ƍo\��7^�v��� <3τ��~�<��Ԗ��<��/׏>������~ ��s�����o��_��{ǅ�=;�9Ѯ�f=3aB�J�Z��ȧ\M��qg�Uӹ瞝�y�O�Nj�z�;����1�+���;��E ׵uFZ�HqcqAa����袟;� �Ɓ�c�0��U�ݠ'�iGaY���+��޸V8���; ���s�L��zǮ���A��G$t!2aT�`��?�Êڃ	S�)F�X�~�b�c9�,�XO��9�- ��}�ss��f��}��)�xM����jM��R� ��sb��A��#�0@�����e���}����"��������9�������3E���6����M�ް� <vˍ��ٶ��T�M�R+U��t�R%͕ʩ^kͭ\�O�cOx���1_��Mu����~��'/�}�'w�󋝙ݏK�4�棭z��]�N%�����t˖�R�\J/;���'��͹41�l> �  ��y��0�;@d�<"F�v�^d]	�h���^l'�W�2�8����K�,aP>�r�atb\�Q�4T���L���Cd�����!0���EX.@';Q��B˄s��b_���= as���xG ƞG�Y�����߂�e3l,��`ɮ/l �m�`	pAg��F�oT�+%6Wͩ�82Yȹ6�AqQ�����0��*):!�)N�.��/��{�֕OH4�8@��AC? ��c��{�ڻ�]�����N���V7�D�r'uj���Z��}ԉ�j�#�����q)*e�56m*�X{�s��|�-�����R�������ިݚaX0Ӫc���'�����87����f�����w�`x��4��|\DA��ȋ���p#iB�<���X`Gh Lg�?/u��ϻ��������bd�0�1�c��t5����3 �V8F�c�Ja�_�n��P��.�l@���o��
�r8����w�3��Q^�+�6��K|,@(�.L>��m�u5_�-F���W�qxs�.G(��<�9y��*�%�u�,�n/��A�Xy��+&�)3 N���R�0\l3 c�\����p@Y���i�Ub%�_�u��z��z?�L�+�n����۶]��5}T�<�zk�E���DoM�ԩ�ӞT�4W���1'�oj��?��i�൜�X�cN����s�+�����s{�����i�*��ޖ�r�������4��ؖ���ү��/�S~�������T��r�8p=�d#b"K�E�sa$�0l#f����0��lh��ha4*߹-����u�`	�8@P$J]�w���N�ŉ�~Unǖ���Z'/�R�	��9�C��d��T^B0���vڼy���/ �<Y�-��}�M�CzDX1vc��h�zbf5�q��=����a�������zl[%.]Xo��)#�xõ���ye����9 ��C<��;����q�xe�{��>Pd���6�&�LD䏃L|�Ŵ��F/�߽�D�����eC@��0�,�T� �ϲ;o�t����hͮ�g2��[ޭ���RJ�R'ͥj�WW�gc�1�8��{Ձmq?�2����o�8�z�֋V��E+ZӵJ��ʬSn��'���c���.u���8:�Fz�ǥ��n��f����Ra!�(3���� \ԋl@����߲#����1)��VL�=��8 j�"���� � �	#IP&�W4�Q@�q�Ƽ����c*up>L���fۑ������(�Q-h�HGqr�g��mڴ)�2���d¸� :� ��&�8��.S.z'�_��O�m�Uk~�{�.n��GD Ҵ#�y�l��[d�܇Հ���p��v��l`㑈p=nX���_"�������m�6('�}'!x,���(C�] s*�͛7�aɶ7z���;jj��oZ����Z՘>�S�)Gnj�rj |��4��33�������cW���\p�(F��c�������<�����wl��W5�{��TO9�|��:�	�%n/U���N'M��R�>�M��jtݤ6�]@Ɛ^��e����Fo'���0V/��wq�.v נ/��	�zq��� �!U�%h�<#:�0&A�c�dγ��I
�B��Aw�ו>��;���#�At.�lLP���>�腗���W�` ������h��!u�{n� ����Ł3���A5�Y�0n��,�d�X~���|t%\tã�CS�y��(\5ʻ�2�z0�D&\x�eH 1"����A62*Sv���>�<�F��\�h=t~��>pRe�7��s��Ww�M��Z�]�r�L��f��j*�}|���Tk;��]�͹G�'�=��;^��~^w]�7l��t�g�߽������_&K�&�i�!�d�x�>�l��Ff�,��Ɲ�q��1�9�>�H�+��ҹ�4�� �я�c�, �L�bXLܙ~���\����OC;�w�S�I�{�b�5v�CY���Z�r �&��:z4����;c�A�:�SP� laYx&HD֓��^H�_�3:VoF�6����w�!^#�Ɂ*��L�+tRz��XV �]H��9Q��F��
�Q��Y�{�6{�a���8���$[��/���x�ٜ��� N��%�����_���-7�κ�;^��5s<q©=;�0aA�=�J�r�-�Ӯ��={V��������>��k[�,����������2q����w�󧦧?ٜ��`���"W(;� ��w��<Jw�	�J7�%��l1�Wt��_�A0C��E�l)�1׈/��|3^��b����͡;6;	D�0 �s�j.�'���)2�����s2��[1Z�/����f��p2v�A���k�J�  �IDATtQ�!u����"��4�5f{��V�c�@l�5��kjkʆ 0�a둡GV�5�������`��s,:=K��đW /�d��=)c������%K����ౝ��^���m/\՜9�]�M�v=U�K��.WR�Y��N���s�D��k�jc����������f�66$�tC��M�R@v�"�&2J?ը��q*hq��GU�6?Z	!T�(M?�&�*�
��T�U�4���!�/0^���̽��9羳g��ݵw�����̽�|��9�y��u�4SH�^���]s���6�۾Y��\ɩ���_o럟8�.^xP�_��?����u��8���BKA �q�тf,;+��t�@|Ǫc$a�lȓDH�C1P� �������Z�� L�<���!#)��]k�׆.=�	�9b�G�y��#w ������Z�C��]�����[�TSDK��-��3��N	���#�7���I��[�:�A�.��~��F>(����o+�F~DŭF_�lJ ��?�j�C���<=|5�Cz�vp���P�����B	=8�SY��5�[3I��v���g���?�	�<cn��+[��=����:ώ6ϸ��P3Ƚ��6�`:����,��@��\ԛ�zN��ު���,����G�vKc�TV����f�>M\z�M|tW�^�� �c��u����C&)؂k
�v&o	[��XNF`R@��gu@�5�_��MGd���I�A���݈ &�x�� �6M� ���@���D-4R6�H4C�Ǯ~�^��	�A�a4B��$)�r4�$��E��o�k*�@G�^}�U����y�\k �A�W� �)@���I/�2�w�JI��m��,=P� o�7�s�<2r#�����>�.�G|	���0ʄ'���pA;F:=�oS��	!&�'���?ڷo��o�Z��Ov杧�?����3�^e�Yd����M�1%{�g�����3�gU�����~�7��w�wYe�_�rx6)�LM�p��or����1�llL�f���]��ӫ��z��LN�U����hvz4Lj�%�0$,��L'��T�I��'�� `��I���#�`R3I�؊��.�`�F�du�����#�L2�0|a����(Y��?���э�ɠh��&�FPG���b��cF9�� -� �>�`���/�0��� ��$y�-�݂W���n�s��'�A;��yi�`�A:a���6����3�`��Z�.�v�$�?��0<S���;T���qz9vA�3 c3�%�K�w-���������_�+��:K�0��d�G�qݹs��W����\$y�z`��;	$O�m�Hpɐ�A&��ix��sΦ�d�R)�a��
�t}���I9<���=�K1d����?���ĮQ��j�M�PZ�F�R�ګ5ZĪjU��Ԫ��R�����V5�ؔ�����γ�z�s�3]��p��i��L�0�zo�y)@TYfvf��LS"-zDm�0z�EJ�Ę�y0P^�3�����=s�C["	��sPD8#���ﾶ�|B�����o��'	w��
�	.�S�<r�qҟ!��&�Rf?i��	��\�Y�N�mO�	$v��ģ�bHj���qE�ʉX�T�($E~���8�kq��~��s��~��VǈQY0�<��wm�3n�*e(��!2Xp)W(^FYȏ�M���ڐ0z��(���1%��Zp�À&�N�[���U�rZ��1�Y-E����X�:�%����Aio��ޘc&��g�����w?Ek��8�-�6[����j�1����?6ٞjW+E��M��q�F�I�6���F2�����D�< ��D?��������+)��n8E�	*�������V�m*����2/��}���$Q�� �+!���6h�I�5?E,�qI�Ʊ�6�:e���� Ì䠀u.n(=�f.oZ�*��ڌ��tZ�O��.x�*uS�ʩdKҔx+��$��ðc����:�ԸK�,��M� \����5(��k����wh�l��h�m��"�Κ-�Sڱ/�G�,{}!����;�~���T]��q��\���o�X!rB�:A~AǮ�w�ґ~k�D�"%ᭉl�4Ց[�<����3�XGP���:��[<��|^�8;�0�&g�7�K��8��B�w�n���aEߝey>�o4��v��%��4D�e�~Ʊ��?Ӿ�CM�5y��w�k�3�����d��%�G�o�=d�;���I��<�G N���v��<������0n�S����'� j���"�C~�Ñϓ(�<�+m�z���{@I���pY��9�qʇ
�#��O|n!�}�T"[��*yy�Z3�g�f�
����<��>�!Y�CF�����&Gk�sX�yy-®����2vW?-�ʁ����g���,x/F0��H��"Ax�Qu�����?�R-��p[�<���1�\�Քۡn�G�f�d�%���{�𞙅aF i��qee��#7� ��3��׏7���;$��iX�z}:��`�����LuB��?���<��("���y_���[9��ED��\�P��Q_!H���I���B-���M�B3jf�={�F,�7j�I�6	)�8�_V����>[����wkZiͨ+D3#�0��0���o��?��y�Ʃ7����?�?�:�>_��~�����Wn�J$����-�y�w-�U�!7�=�K���62���U�f��7	���	��I|���*,-�\eF�I�G��Q��x�銃� ���}�tW�B�� я�<�.s�վԣZ0y;�pE1��±G]�x~�s��duF1�T7�N\P�����K*�d�5H5��{���៏�d'O>���͎���xr�&�{�կ�B�;]Iwȷ�*{���Nŭ? Ѧ�Y�6���5Ɩ���Z�g�n�M���d��������̈́�+���]�&Fܣ3��ȝ����\��m�����J%�7�N.V^���lOI�W`��Ԛ�;��rFM�hO��&kSkwK�F�d*�=���e�yU�2J�~��s�<�<�m$�ȁb��A����F�1$�JCzG�9�0�X��=@��L\j��nl�˓�7��d��4�̈́���=E@���Y�����Y_ވ�o��N?�vҖ#b	�
�{�� %�R�o�l��u�i3����7�( �0_#G����W:�z�F�I�Sh�_���Ĵ-k	y�E����uh|�wrn�I���K]���+ԥU)�~��J�M��h:��,���0XyO0a��W�m����m�	i[p��������b�w,wk�n�i���2���|Q�aӿcOd�����ޟܟaP[_�BV!�,��
���I��ʠ�5W� �>���O1*��T��C�".C��±�$��&�^�o,k���`>������b�=`"���r�ʼ�"���T����n��րj�����B�������!�������Ѧ���C����I�ǯ���>ZHc�K�V��
�;	�`"���X
���/�����$�Ďv,�[��5�8��f!�-F�[i^�G��b�#�ۣBb?B�/_ɋݭК�Gb��xI�ݩ+��@0Z0c��]X�)��"����lps�lU֩ʑV
�&,��焾��;�E��sx�g�k���=���qH��/z	B�=���@�!7l���������Y��K��WCNC]�����:�0�w��0����ɻ	�%�e�4��()��c��+iY��l!{8� �j���%�&�Z0��ә�<���Pf��36?�[�z0�M�?���x~[�੓I[*�" ���.�$z��Y��f!1����>�g���D��UgΔ��2%z_�ֹ�\
���82�~Mg�kTZo�%s1�ˑ������ݣNw-��)k1��o�Z�F&WК����D���i�5j��W���r�mEwm;�u�`��IP����P㕗~��Ka����B0�A�q&�>B.���0בTI4K�� �i�?�R��1u�03<ԏX�7�˂%'�mj�9h���^����ivJ��A�P�4R�m^���P�MݸY��� 	3�ܩ��^	���E1�5� ��$q��lJ�O_&64��%*�����b���G��O�w��;�����F8P��cfpBiN�-1R<0#-p"ϲ���R��,���a�F��IO�sd���e3����I�F�]&�N��74}$x{L��*۸9��ԃsNVق>����{6�k�9�2���[չ��y�0�H�e�UKGd�V�)��
�?�R�:���l���<XIZ����l�j����A�h���r�W��y�8�X�;��쎈~�)S�v�O!��ێ}. �B���t&�Y��)zG�A�2y�Ÿ�3y�`�
��PeuW��.�id�sĻ���r������!?j�6�#ي�V��}�;�v��#7� �eqe=��q-MgDbc�,����<�=��]79r˫2���x3�ȧP=���}���u#AQ+��|��CQ}�Qűq�E���Ȳ� V.Y`�F4���w��o��{@���x>��	t�@h��;KmO+K�ҷR+��6,.��+2c��A����-r	��Y�����WZ,c�����2�*���1ۤJp�����h�J�������Z@�8�/ILM�����W�#�'�����J�|����q��ٱtǀ���Ϸ9��wW�wB�B�lk?%���������Κ�ꨭ5 �_R�F��Ԯ}�3�"��'?�2�S�t���(>����Ν�O��\��p2Z����4h~{{��8Z>��#@�Πu�Π�S0�.���sF	Pԭ��d��H��=��PX��x�v��o9q���="�J��[P����{ǭ����;o���NՄ�6��.��mE�������Ҩ(���<�պ�?	~�W�-e-6.�$���ɋFaZZ���?Ǜ������cU���!r��鐵�����ʗ;^';0i9fI���i=XI��ɝ���:��^�\�n�{7��>Ԋk�����>�;��Z_���0�7(penHV�3�Sx:�Ҹo�<��{@A�4�t,r�A���hqb�&�au=��S��
��.��E!��;\�(l
R�Tݖ�V�^�h����Qt{J�~aulM1��Z�'�}��:��~ϝz���I��`�ϊ<O�.��GS�؜��i���{�k��	�;�j���\�Դڹ�,`��>}M�=;?֘����D�bZ��"��V�aH=��ov��,w�pn�ө�o�Q�+�/?$U䴐�^��g�:ںf�c�j��д^�w'2�_�&.F�m8�z=E�T��|�����^�*`���r��.H|):�F0�ޟ��_�2���2B;���P�D�	��3�'y̭]]CGmIR�����B�|v^�=�}	�߯��5��M}�XI���n���2�S��ToO����ޖ��_E����KPɸ����Im���ˊp���D�l�"G�,cC_���G���)��ui|ۯ�u4�Q@N��)j��3�7zœu
���hPۋ������|�q-#&�1E�vK��/j�ET
#���A멃�,*-^�!��GA��T*u�*��+�6�6PŁ���\e4�Ҕd���x益�������m��Bj"�7.��̗m71�!��U����;<��o�]�K˰�u������������񏯣�S��FB��tC�_WW/鳇Z_� Ps��k�Ѝ��x �����ö�nv@9��s.ƒ�d�������%��V�C"��Y��n�qX�6�G�?��n���$>�z�c��,� �WF�.��}1�{����
W�+g�VK�Kb��6����w:Z�%�Ko\(�[�s���������2��=��($T���.q��hB�@3%��]d��a~~GIɿ$�Y����������k�*�[?Ceg�3��rƔ2��v���ގTڵ`�M�oOl��PK   O��X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   O��X'�Sz�  m  /   images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.png�WWP�E �$�.��(U��TAz/�J�.AzI(FRT:"A@� ����P�j�b@�����>���93;g��즚�2�x@  �Y_O�좺_���"�\� ^`��m p����ma~r�ޱ	5�E�{ P(����o��K��L@���-u �対�-��|r0�����|{22SԈm�����J0��d�]��r�2�~�:>������OT��9tW���,&Z��IB)����Me�iQﭹ/��G�����vѩ�6J	{NԜ��O��:(s$|�T��a�k�W�jjn�cX��e�!|�1��/><=�Q�����uu	Z��y˜��{����Z�xc��8ЮP!�Pݏ����]��J�x�nUz��tY�KD[N/�!�n!h�t�-�)�ZT����HXQھb���3f����cn��r��:����?L����m�?����#"�_B>������+ń�N�O�	'�a�!S̡�ɳ.?�K�+糮_�1zU.D��R��s��LM>������IZ�Uy��N�ʻZ�=^1����&��/�j�{~�B�6�$.��h�	b���K�
�Nv�5<�5U:�ش��ґ��]|dӏ`U�]g9N+`��&\g#�&0Ii�~Wi��qF��G��Z�ɻ�<��=F#P��{�q �?�(/M�fś��&����ؖ@��9�C�L�r�KV�%���gV3)"�r���9���A�1��K����&�̑~G�ZS��`����z�@������2\c�)��u���fY�U���J��������t����N§��r��n�DT�ם��I�4ca{�4�R�/g^�Z΀����*�]����6��H����4�����ђchw�n��In�9�6s�kž���s�_�q*�8lJl�$�B��J�^!���g��YGTW��{�Y�Kv@�~C��N��p������:F�I$�y/���=��}e���!7	a�y_�,D!����\~��G���1K���۽��P�1�^���K��]/��gi:)/DT��ձ�W��4�e�����׻�TP���N�Ĵ�{�|�~+� ȿ��TfT��_v�]z6\4�^�(�/�?+r�^�-�R\+�d�߮��`vͫ��I����R�2���#�:���\���/����2~�ޞ�6�OT��A+��U4 �{��V�n�L�9]	&u�Ê�ʁq�c�IW7F���&�ڿ����:�}؆��٣��C�ܚԟ[k�&��>4/irƛ#r;���?��!�:�Q�n��j��p<�@B�0�?��`tty�j��~�✫~����]�͡����}�`洴z�hw�S@'2f  ��!=�7��r�\�pW�쨏����C�����xI�����TIΨ���Q
B��������������D٘!��|�^���t/v��_��M�����-9
�ںmE�m�K�
��{�(��yw��2'�y�4)K�	�WN�4{~G�"��p�^T��W��z\O�g�Җ��N��?��g�g�a6j������o{��xq�VD���r<Q�R�.Fw�����X5�͑�wQ�d�@�ݕ�0(�!`�5�6�8�.HלI96�<��X*����AoV��W_������ɼ|����.$��ڎi���J��Σ��j?��1��Ս��tƛ�|�;N1b��3c	e�~ͭ�W3ɾ9�2	4�';+�~1?מ�\np�E���@�9���4��V	b[>tҗ�Ψ�\n�O�G���B�$�ܯ��l����bH���r�(kDJ��o��������50qu%�Q&�l��q
ah��B$@��T�>3�=�KR�a|D,�'�RD�7[w��p�e�	m�`#6�-�z��/�R��I�A�S�ݥ6������H�G������׸�<Ի�}͒A��)��?iS'۹�dq�@0�p���s�uD�EJ�~=��[����\���Ű�˺U�Q�>�N=�)ߡ��h����Q�C�t�V�g4���5".TkN�l[���?`�z �"�����9�� ;41�r�0Zv��͝�9��E����hth��kK��iea�a'v�/IT����"�R�aQ�2��Z7�M�(�@�8qf<	҉x;W�+�\l����?��߫�å��^-MW��<������:�[��(�Q���h��6@�2zP]A<,��3���F��[��~��6͂�J>
өQ�Лw��z����	8��/���M�W�n�=�ѩ鮎(�O��N���'�bSK���%��C�L��M*sޞ�嚖?Js6�.Hz#�o`�]�k��Ӑ�J�}�gA������N��[��j�
���&�u�Z���,4K�:&��V����W�����w����'dӧT(��ϏvpI�1"���ԥ�[�N�C����l^!����d��[N�\�������y7�s�������!/�B�'S筱d��(
�f�Lc�� �ϕVG�֜�y����Y�W=X���C=O�x�?�}�Ͼ�T8Ab���'�r�}����+n����o�8�n���Q�8M�ubC��S-Wׇ��Y�Y�^h��K�[���y'�>0B

�U�d��� �.Eo���v�[W���
��mYe��>=Gc�ְ�36ꍽ�J=�U1eR�ѲoR5�q�DL���>.o�ps���t��&�V$�P���s��H�3s����t���kJw�Ɠ �K��YK'}4�����N�; n������`��~�Py��S>�_}�ff���{-��h�YwaPg���UAt����#�c@A�τA�5G`��{� �'an�')�,�8��&���2�>*BaW�c�C�t�5�0m�niz���M�c��I�0+�Ԭ֢7��q��H��d;�s�~��q� ������83�{�h/�#��nC��H�߳���v��M.�����l�ýM����,{�	�!b:@��LN`�gIZ�I���]�MK��͚o�/ܨu?�Sj��Wbo�	���ԠJ�1/f�S|����ۆ����VL�
��d'�ߩ�y��
��:n�P&)����fb ����T��>�W�Ŋp�/��>��R긥��O�9���W�J�W;�Nff��^8%�Ƿ��R%Ґ��&�YBi��3����a�����r{t?�)��⺜�D>��avN9��/:G�
]���i�alMzy唣���>2=v��"�DD����MG8�IYfڑ@:��?X�:��[t�<�MT��h�v#�lk�.��k��j�i79N�n-N�Չ@�ۇ��%
���!ˇ��&�M�i`,���/���;q�t�쩉�%��v���^���`5��o�½���gnΓ���W��������5������+ŗ#S�k�#�g,=(�.o��?~�8�~PdbM��z�S�Q���i�v�o�ք#���Y|�n���xSS)P��Kq�1��J0D����[Z��u`��Gmo�$}�:����8	y�;���7{�?Lg�w[��w������__��;�1A���M|��gJ$[ܣ��w��{��M��&�-VL�FB@�L������5��_/D��{9�|e��\�s�i|mx�S��9i��X�z���R��%�sہ� �1�l�]��5�^� ����ɲ�5Y9�9�M�G�V�׹�{����Yc���7i#���T�S���Ų?�D��^�ˌ{>~�!��82T�;����ਊecС��D�S���W��X��L�/PK   O��X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   O��X!�	2  *-     jsons/user_defined.json�Z�n�8�ï5�/yk붛�M�45X%�������� ��H�]M-����D�C���о�n�Wnz0�m��[�|Q�|:���֛�*�NpB��f��C7Ӄ?n�>��z�/'��n�E���!ӯ�7���ϦEU��C�Z�x���X%c�RʴM��q��UU�r��[�5��;خw�~Is����jۮ�a�'E��ʈf�#�Q��2���\c��MV��+��l'Q�Q�r���X���rE��^*p7��^�O<{˿���2�}wpwU�����7�rw9/6���~[-!�S�Śh�pﴺjh!p�}W?v�T�a�e�.��N=��5��bY?/�	�5c�%�]�)6���{���w�[���؂M�^�'xN����.7��?�{�i _���?ßы����O{�y ^a�{�E ^G�޿|�7��?� >�82��oW񍊔��%0!bx$���Wȿ��HP���0a�D��3�LLx$�Y�!dc""�_�$�d"���kf9���Q?~��rp�'��]3��/yX��r�L�?�����#���g#���|�,b	�EJ�V�����(�:����@��>~�Ǳ���]ˇ�RD�~�����n�%J�$2>$ ���E_����'�aN���f4�]B:o�곶�*��R��K�j��ۢ�q��E<ms>Q��&��j[�'���.�Y�s�ۮvۺ�yү�.�m�r�Y��Z�%�"\���O;�s�L#���T+�#LS���:�����j/��47�a��#/$47uod���(,�W��&��l_db�����������9�I���ӽ=?��\�D`դ��^ ?`�><�\q=#
B@�كO�b@�"8I������͖���x,��_|7W��g1؈�ʖ(.������n�|� 5N��nʖ=�	��/t-�lR���' �@�^���O��NF�D���f��$:��0�M��Q�뗢����ӽ`jސ=�$P����4������r������6TBD3�Ե7!�l à��ЖA�����wm� �@��������D��7wǡ����v�\����]��O��C�q�X��v_�^]�o���={],�M�.������k��}�~�>F[�Ͷ�uSd�S�?��j���{ZC�ݢ�*M�'�]�U�U��>���L.�ZZ���@����?���H�eL9ϐ:C$s��(B�t3�%���:�"��G<K)�;Din�ɩ�\Q��qS]v��Է��Y-��BH�g
��?-v ~2����.�L>�-����&���)��od���+�����_c��:���+Ġ\��(�A��Y���P��6:lt���a��F��6:�?qا��	� ����:p�SS�TW����j�1��e��$(74Wa��p�Ng\��XC���1M5�a�}�Q*-J���z��C1�(��(]���3��P���Z�������ȧ�BC~!�Z��J��f�	᫸/$k�S*!�9��8HW�"+�A)�ԑT����'���Q[��Fm���5jk�֭���PK   O��X���  պ             ��    cirkitFile.jsonPK   O��X ���s� �� /           ��  images/25c207d7-bd9a-49b1-b471-35e2df67a92a.pngPK   O��Xs!��}  {�  /           ���� images/330d02b8-4530-4fd4-b6ae-26fc03cafecf.pngPK   O��X����(w  +�  /           ��U images/42266fcd-641e-4cfa-a619-b442e1b7bf10.pngPK   O��X+���  D�  /           ��{� images/5cebb09a-e86f-4cb2-800e-22da09d26481.pngPK   O��X��"�IY eY /           ���U images/97c183e4-4c27-495c-949d-3fd800d1ff32.pngPK   O��X`$} [ /           ��L� images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK   O��X'�Sz�  m  /           ���, images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.pngPK   O��X�+�s;  z;  /           ���; images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK   O��X!�	2  *-             ���w jsons/user_defined.jsonPK    
 
 j  '~   