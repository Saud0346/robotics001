PK   7��X�����  �%    cirkitFile.json���6��������z�7��6�7�e3H�܇�AC*����3��?R~I�h���݃C���b��OŇJ���*����r��?��z�\Ln��N���S�NM�����~���m�?���~'�?\R.?<,n����VYZ�$-E�ȊgIQ�21,/�)3'��>�ܾօ��Ug<�¹�:e���,ϸ�e���>�h)ZJ�U�)2��47IQ�,1eaU.�E텇���0V��,�˪Ly��җlj��Bꤐ%Ӫ��ʙ,T�,�Ʊ~�CDc�F"�(9��@F�K��k���C�{"a� a�U�
�ڡ��'�q�'._����i��u�d^��VV':cE"-�F��Dԩ)�ҥ�ʷ7�d�)9:JCJ�8L2�#�}Đ�C>d��1��WHy��7Hy$~�G�Ǳ>�G�Ǒ�q$�G�Ǒ�q$ɟ@�'��$5�H1���3��xLѱ�p��)5�`������Q,�|P%�A�����)����`eG�S@ec�!�J"(��$r���J"�WH�r�R�J!�SH��?��O!�SH��?��O#��H�4�?��O#��H�4�?��O#�3H��?��� �3H��?��� �3H��?���"��H�,�?�������BT\&��"�2S~�[�ri���ʣokTV3md�(Q�DfE���IY�˼�m���`��iwd��:�^bu�E�����\�V;
Qr����=\�RWV��2��yY%�Y�;�������x�m�Y�e%,5����IQ�E�Ve��B��1_�U��X{����{�l�a���(9�^��.�@^�l����*9������5aw�%�EbO��emx�3�����lJ[X��s�*^yH�Pg�,����cO3��%���,��%���,�:��z"�R�x|>
�P[�8��E0i�������Ư ��1e�t�S6ʭHj��~9�lT	�y5�r� Pɱ�KV:��Im�Mdʼ+-�L
WW�w�3���т	#��h���O��3��L���'6=B柫/M�!��\Η+dh����2ǅ&-�?��,��k�F�[T-2���5�Ȟ�4�u�M��)&4�b��q��k�	��04�@'�"H�H��U$�h-&h�Tj$�F�Ė��:"xi�e4�2~��QCC0�A�543�9Ŝ��P�i(�4s�9Ŝ�bNC1��X�P,h(DS	���8��Fx��}��5�O����A��
�Q�P�[\�54K�����Q�P\r[f5Fь��K_,i|���Œ�K�Ŋ�+_�h(V4+�Ŋ�bEC���X�P�i(�4k�5Śh��bMC���X�Plh(64�ņ�bCC�!�f����Plh(�4[�-Ŗ�bKC��H14��@K�Oc)��� @^x�f<o40�-�@��7�K�4��;o4�-Ѐ���;_#h����!�\|��Ad�ߖ@�l�$=}q\��khiF��(#Q�5�f���b�0k��1p���1p���-(p���-(p���������؊J�^��t���nʳ*Ҽ��-��~�q-�M�qظ��{ܬ�92���_��k�k�X#p\�Y-����5ǵ��ih\^�e�q-x-�D�$ѢH�h-�D�%ђ�PG/��_F�/����hf43�Ŝ�bN�i(�4s�9Ŝ�bNC1����P,h(4��ł�bAC���X�P,h(4K�%Œ�bI4#��X�P,i(�4K�%Ŋ�bEC���X�P��v4+�Ŋ�bEC���X�P�i(�4k�5��Ś�bMC�����Plh(64�ņ�bC��FC�����Pli(�4[�-Ŗ�b{�bp\^��7и������Z�Z.��k�k�h8���Ɩ��58����C�k�k�80��Z�Z.K��ॡ���x\��/���ǵ�U�k�k�<	�Ƶ�\Fׂ�Ҷ���_��ٞ�r?����r6�|�����a�����-ʭ&�o�:�sc�+��^DJ������^�k��lA�?�TU�B�4�h�5�8_���C<1K�H���9f:�)��3�=j�):WA��C�-q/�Pec���6>�����k����5���)9�1Wg�23�Ĕq'��A�d�3���\�`� ��3pDgd�~�b���ߗ'_n ��Q������8�Ut��������ݕ����׻��Z���F����](<f�s,�����<Ǣ�ص1�	�Kd<ؕ��6x��Y�c�|ր�X>�8���?�ϲ�>k��	L�.�	L����'r�}5� ]_�?@���OG B ��[Hr;�jqT�D�� � ��y�a��ϱc��Wc ����#���j��&��M�{��]���y69�6G��g�������,�p���n�v�a�>X_f���0?�2P��|���0`���q�-���c�*>%VY�q�y���Hy����ͩ��1���m���髋L}�Gg`�>ò��K/��˰�6a�(
�@c�,�K"ǒ��~K"ǒȱ$r,�K"ǒȱ$r,�K���(�C:�D10��~8e`TGmb����t~rŉ>�/���<�:��B-����j~�ŉ>�z�u��|%��J��X�+��*,�
�|��*,�
K���$*,�
K���$j,�K�ƒ��$j,�K�ƒ��$j,�K���h�$,�K���h�$,�K���h�$Z,�K�Œh�$�3$��s8Y�D޼�v8Q�� �� �|��:�'�"��8Q���|�:��� |RDW[,L|dĉ����u���N�����n
ƺ3�@	�|�ol�K�>���)����D�`h8 ?&P���m�O���/�H�u�>��D]�O�� T7`]lP�[A�n�:�8��U!���_�PHd����$<����a��D*� �ˮ�t��_h��������h��Yl�f�lXm����ǡ�Q<H�Fw��A�	$x��A�	$D�AB4�	$D�A�	�A��Y�槤d��AB652H� !��2H� ���
*H���AB	$T�PAB	$t��AB	ݴS��AB	$L�0A�	$L�0A�4M$L�0A�	$l��A�	>�@&���� ����# �Uv ��H_&�iv����n� ��%����֍,�&x�{3t�ɿ �� -L$&V
�o�i�Wy��3L8S�x���Ԝ�{�ak�� ��[\ �u���ak0_a�<��_Y#*��
�CЯ��T��fĬ�����ྂ��;�+�ż��U�_���L���s����s�g�cs�����cpߠ!�.T$6j=˱7�ͅac��$���+�Wa���1a�E�	.�-H�9؏��k�M8ct�n�R�ɿ���n�*@zr��n��-��������ߒ�[�K�n��-��������߲�[�+���z�ؾ5X�9ء9�����������-��-��M��M��m��m�������������������/<;�|~_�\^�|�⩗���z�]���H]�o�s��f�|p��̅M��{���l3[.|ƴ�a�d����A7��ɖ���+oV�*�.�NLU�e�%7V%�I%���U�F:���[��l:�-֛|Qn�v#���j��['��o�7A�lU�ݮZoY*̍7��驪?$�Q�?�
_�y��g�_6��ly�l�n�M�9�>MO�Pb�J:���Nk��aG����ʴ[K��:���nkYu���?�j-i�M����R����=񴖜|xX�����9כ�l�7n������|���{Sh�1����'�j�~���w^����k�o�����zV��!m���8[9�h�գ���!_<�y�y\�Ӿ����,�~IK`I%�2�{�4����Y���,�D�)Β���tc��<9�A^>�����E�<�T�x�[鶕��;�+�J��tӺ��<:=�k�J�t�J׭tsL7i��V�L�^�U/Ӫ�i�˶�ͳ�=[�ݵj����ֆ�uzL��1}k��Z��E+k����m�M+]��e+���wf�ki��Ҵ�U+]��y+��=��k{L�~�<^�V�n��V�h�����;iڹ�w�=��K�V�l��V:;���Ɩõn��V���M��꼽6�t�J��t�J����P��;�:o��Q׮��k�J�tvL��y{m[麕�Z�b;CYV��z�7���ʭ����{7����w����dz7�UMJfLb�D�ү�\ʻ�*��J�J�M����0_zo�_���;Y�
#+�Ty.��T+?L�4)�J�q�d�l(�%'k[�:�aG�/��PI^e"a�w�u!��A����q�֜��]��TꅍH
ckozZ0旼�˶\�^�삊}����cM�{?�W-͵�d^�<a��f9e��<1"UU��T�4�w�j������F�4ϋ�%��~�P��LXߴ���T�c6��|7_�]ۚ,�"+�4ɝ���"͒L���V������rW���/*�����v'R|��?��X4w�������[�H�s�s�I�Λ�j���Z��zw�˔j��l���Bm�|�rcs��<%&-a���)!��M��
��ZG���D�ڋ�~6�B��g����K�e�yH2�|ӗ�������8oJ������b�S?�³�p`+�ϥ��K�\�'���y7���U��n����������ի���/�՟����Ϋ���{�r�W�������O+n}n��/��4���尞�l1�f�\�q��϶��忸�+73��_��t�u����&O�e7Y����?���E�q�K�Ly�W��� ���QZH��eEvÕ<�LR�(�qaŦl���eIU�'��f��2�$T���f2d�T�	�$�֧?\j�����q
�1Cp��"W@F@d;��"bҿ���PGD��>@S 6x�fb�\��#���O��B�ċ��b��܍�S#�J
(T@�v�!;�:���8r��7��]���~��_5����Xnȡ�}�o2��ݵ��~���$�S�M�mzL���O�e�<�:�]W��:#�p5�P��)=sW�7_�[y��^���Fji8��;��{b8ϲ]��l*Syc,���mZ$�0��H�=�6M�H>ioK�jv����ϵ�����w���*��1���d��w&g��&���f�TX~cL��ސV>��N���Z����uٍ'���lX���5~�r�k?�<d���M�dV�}�{m~�+SgKm~��i?WmB.�v����V���2�(�J�-�_M��!�/�wqFz��Z}����AU��0͒*���~�m��'��Ζ�d�r�GFp�~��@o�����]ɮcms�&J�����򶉶���
>h�,k��R�f2���u����z;���!�Gl���	MZ�j���{�������c�$���wE�.�Q|����擉O�j�>h0�	��i>�x�7>�s}��¼��S�?;��w6y��U�޿�Y����_g������	'��^�|�j6��)X��f�7�j�f��mY=9r~��Ϊ��7�V��_(M���Ag��r�ؼ�7�]����&!���M��K3�Z��۷����`Ӂ{aۛ�!�t�-}J6?�g���r7��B�1��.��R�8�.�1�:$���z7��ąl_��ח�c�uׂ�$�m�y�ּ�������'T��`ă
#��dPQ����'��FŽF/��^��}Uh41�;���	��
_
��]�^�a��D���P�,sF�FJ����l��l��F�������t`.��\�x�ѹl)S�N�J�kZ��'A�ۨF��)5!��:j:���ၧ��\���?�g�O�外�i�Y-��$��a��}α������*�R����x�� ��p�F��@p�F�ӊ#
�Ԋiwf+�d8��ՙ�	^�3GXw��l���LX��KZ�
��痺����Fwy��Z=8�4�\_Wg¾�}��a�U:�B�}~s��i�r��&�.�w����|�u#������w�L�u��\bp�
����u~���>��2>#L�3º��t��AHY�ts��"� ;H��c��G�F�1�4���ªy2���/ �ʆ���LX��y��#�a�'x��Ũ'��aq	�X���P�]�_wC�����ξ�ݾ��l\�!2���'yr���\�Mߘ\��`B0,5����˻ݩN��!������3���%]�K�� ���.�4�v�!��3�k�?hu:(��Knˬ&�tذ<����P����םg�9���\�N�\s�頓鶉�t9�4�m�'u�!�z�N;�^w;�=i�:~b�]QÙ�k �a�[{�?º��N/?�:y�Ӊ2�dʆ��L���m�P��R��3�I�/��뮁�݅(�6�[�͙Z�s�������r�F,���%��p�Ǝ]�NzsT�� w��+6bF֭VT�:��n�7�j{'�'ѡ�$�e\�>��#��Q��H(�#����.���6�N�����A��a`�L:<��'�=�����ke����SF���I��÷������q���΂��'���(���7	W�ug�.�3������c.�[�#2ۅ�KN?Ӗ��m�l>���1߸�,��'��u���߮�1_<��o�^o܇p���w����]��ޭ���a�!����PK   7��Xs!��}  {�  /   images/330d02b8-4530-4fd4-b6ae-26fc03cafecf.png�g\SY�>�cAQ��� *"�Q�Q�t�ё"�"B��HG�N���'�(�.%DB�HhI !�?fFt�y������0�!᜽�^�Z�j{�]������^�n�����[�%�n���-��ߘ��I��z�73�u�,/����:��n�Ⱥ��Ս|'zJM�~�K���?t_F�a�ŝ6��<�x������ޡKw�Y����֡�i��WOt��O��3uF�.�?Jh;�@>Y��_�#�5?A��ۙ䖥�R�L9ɞ�*�4�?��Y���ﾫ��o��Wm¥nL�n�k�R[�a���u?�qxS��ҝ����RR�T�"�n�����oFio���?�q�٨�S������ׯS?���Ư�[��Е?�)QAcek��h�o&��쏮yAH���;_ߙ��N7!ѹ�/�m�߻�����3�ֈB٘�<��%�j�7f }�KZ
~~,ۣ��ˋ)ybz������N� �e��A'���ˣ��.oH���f���ʞ4xd$�U�<�o�z�1���ڵwS�9a����8z���J�2���y�u�o�Pyz`� ��b��*o�G�D۳��/ep�cҘ�ܮ�%=W
��c��T��,s��;���#��S�'�4��,�)���\�jR�zK%�p+��5�'x���U��u�G�Z#����>���ԇ
^�x�6<H{��v����"�䫇�Ed��U�+'B��"�����3���O�7�65�_��E����1nZ-Z���Uލq�Nm�ě�}�̦�Q9ec\�PsV����퀴^��>l6߿ӦИG3��	�BĘ�����p�����v	��I�Q0غ���6i/Y��&��7��vJ��x\��٭2z}�v��H�?nP�[�#�-�(�'�=z��z&�l6�xh����/�� u.�d��8'��H��/��m�j{���$�E��M��w��A�7��~[���IФO�-w��$�6�^�!<�l~tyu'�i�coB~b��X1��["�c,C��ň1s��x����3�󽿵*�����G,�7]h�4��f��T� m)KA���~&��G�g���U?�����ų[�;m�|�DF��gS�dD��Ŧ<F9E�d��ݢ���J�����홈:y�U�fz4�&���ھ7T��L�1�C�����~�����K���q迪�_�����6��!�H����4+<���F���֢���7��ߪ�)�Ѫ�dSW�.��<��[ ��)�/��;D�[�Yfŏ%}�z���K��:����m��q헊;�����>P�/U�C&<d��]=�!��1wڂR����-�J��Q�r�>d��E6P:�L��^Mu~?�/�|X}�k�'��6ɑ������]��hC_�����o�	�.+ae���v"m[m����5muk���}&�n=bx�c��l�	αck�~R��'��ǇB�G�������1���R�`�_X!8��7�v>̩U�[.�8r=Uz����ȳ�(���Ll
���<�IKj�~L�{vl��|<�k��E"Vcɳߦ������Z�-.���m����k�#S2ڃj� ��ئq��9����6L`۝��/7�͞L��(�0 �R}0�|0�yX<����G��I͕�v�?�Fr�����t�H^�_qLt��{�;]v�q���1"��	N�����=���������1��ú�7;�ffE΀��`�������B�ٻ�1�D�[�kx�:#��� j�/�:/}���PR�c��t� <D`��5�H슛V4_K�������e���0�#mu����Aڼ�	E�H�a�����7������-2ծ�H�?FU�{���
+˹q�ѕ#2���~L���<�S͏����+ �q���?:``�',�:�����{{�Į8!��܏�� �iC���\���©x�//�h_�Twj|�`C����L��OD}^m�z��i+z�z�P���l
���0g���\��Pw#�x�E\> ��E���]qGd�V�=P��+��:�ds�x�䷈1;j`؏�����O/o�����׺Eॶ|t�C��i��ZB E6{�z����πsQ<�C�;��䐘�V��x�����]����g�ͅ�M�iB���=���Pƥ�C��T���B������D�=�=��I~����:���19v� �;��~tL�o��'���B��!Y�k�c�5��WZ�D��f�܇�^^���8�a����YB�b��'�"�?z�s���P!^�IRS��p�t���6�����=g�C��k �`�A���|��%K�����W�����U��*���
�_������>�'��>��"HO�8���}J)��ۗS>���d�]Pv��wl©+���qݓB��zj����:J��$��	��pwQ	�J��S��0B���w���І�-��(.uBſv���"k��=8b��IPZ��s.��m��Z��iyb[b���fޟ2�]#Ž��!�}=D��F���<%D%��Z�xڼ<B���͒�>J똵�����q�ź��e!��ʺ̘�!�o�%��h��9��l]J�������|�"�U�c�\0�D�=�z���&f�a�唖��F#u�eNY@�Mc��~$'z
i| �k�w�Na܁{�1�c���8�r�)>.޽�kcN6���ʡ�wh�_$uL`�����Ylhય��J��X&M
T�,�.�1��־v��}����^�|�B~ν���3|�]KҦ��2�G��n"a�QY��е�G��Ӱ��'D*%�^<KF`}>�]�F^� Ŷ�1��"E��p�K�Ot��A�B֙Z�������a�w����r��\���8��Z����Qd���(_7�/$ת�f�����jQ���D�2ݨ����E-������)Y^Uۙ�B��nٽ�^�Ǌ�pM�H�gG!��5����O�9j������&���·,"�ӕ�j�w��4��z��kGSez����]�X�̠3�I��l��<��W�o��s��!CQSx��Y(������rw��ˬh\E5��Wt��̓��9k0��d _��ײ-Q���xfr.2��/8�� �<����G��?���]�9f��S�-E������6�Z���/���ʶ���h F�(}D&iKpi�g��??Y+������X ����v���s�ٴP��"�ϥ��o?�`/7�l?~�oJM�=b�霤]C��Zu�c��@Wl�B�~d��Ԗ�¿��Kk����F�����h `VХ��gL븖1��:	X{$��6}"���![}��#h��LŎ��#̞�Kk0��?V�=m� ٥�����o^x��I{ǈ̆3TV�����ŏ�Tz �b�iZ)����<��#��\�]sn�/�`K���2�sq�f9��)�+,�c���F^�Q5�=e��!-�[���q2�f�����g}�Pr�)���Lj]H"�л��隶��Yl9�J�����kj��>����Gr�zGg;B?������-�{ײ�3#2S�$h��d�Y[d�<�/+��qԹ��<��Ι��T�O��ħ���ලl�~֕�6KD�}��.����H����Ԭ��w
������e���ǸÛ� ��؉�1���{��pj���{����9���>L���O�8�s�1�)�_% J�R&+�����D�M���þ=��\"+~���Q�r}�Q�v��f�L�e8��:Ǯp�뉟����f��>���c
5N��p�4u%�n(B\�}��g/@:Q�h�`�piu_g�q輡����婬�?*���gG0kx��?�����s{��_�n^�L5t��6�G�N%,ؚ'tr�Ҟ��S=b���@��1��(����F����6(Vc����Y	���F;j��Q�'/T���Dv+yA�v��}^Q�Ӹ\̓�2�)g�\������&�w�����a�1���i�l�ZKA�S�Ez}H��D�,�Hr�W�}O�E2�R�R!W�X:Sm�W^^���N�d|%?�W�S;��*;�Ayt���T�u_eI;�><7P����ɶ�E8��E�iఙ�a��I�D���<~�Į,=�$�p]�=	7�H<�G�5� /^��[Q�u!,�>~�*nљhΜ����{Ո�nz@��s������W�{���GO��H�f.�������G��P�����^j��NA��N)��X�VV4���>U�gf%g���Λ��4t8:s��?�p����c	$�9��6��5t�䰶m&i���^�����i��.��4b��z�P��
���/Hrx��l_�1�\hoEu�t���+5��yh�8ﮖOj䦠�~��ݮM���Ġ�4�8���-���ړV�QPa��L�[�tC'	#K]8�����a9�؟������ج��f�/<X�E��ZbЎ�א)P���1z��9��7"b3��~�?���~��O�)�	3����dØ|RKO顊ThU��kc��=ϊ�e7����8����Ɏ�-�N^V�2Q$�cʕ���w|؇7��*���+��.J�k"<�nDo>�=�Xf�ȟ���g�5�߫�����L��|%���}���D���]���LǓ�P��+�}c�h�ư_l2]O�� �jH�/��y���/u���`r�it,�5�=�`o��
텳x!�[KT�}L`��9�F����f��ڳ������C�/��r��F�#�e��Ļ�w�ڼW�^�'}A~�Qp�=ͩ��U��s��\�����5Qv�����,R�	�2���J�jp���8SLEk ��L��N��k:G����G;��#a;S4�j=Mlw�tﵶ"�MX�=����)�Z�u�a�E��"�`��f��ڵ�EM�#�$�S >p�����)�b�X�-l���^h����q���| �Û��v�&U��(���
�c�h�}��.��`�G�D��d�R��H�l���y��D�����"{�3g!8�YЦYH^��Z��6Jn��>��9��:6��Ά��0"��,�g�bה_om��蔞z({q�U|�\y��n(��P.��m�C�iΦ�Ѿ����$���}�v�{������9��؞T�b�01b��W��N�H�@���B�=Lݩ�����c��I������U�_w'�%7�X ʛ[+|��,SQM&t�/���/��:��>H|�YMҺZz=L�7�fU���
�_�xE�@�<�՗�Hs@�r�)O���/�rq%��*���n�o:�K�����(��W	�J@I��v�:�[*�V��󙈮%�����;��F2����Wo��$Z��B�~�ҵ��NT�h�S��}���#��(��8�dc�T�_�bئ����4A��$�Xs@�Z��/�&�����e��[)0��0��W1��D��[6�:L���s	�ӊNw�;��� ���r�^�%{�Ȃ��]f☷�/��e}�㺯�{�bR��B�J�p�n�;������U��, �ژm��1�a��ܛB��!��UU���e¸�Z�]�����粧��,HV*�$��e�y�6a&?�1�>�?�N�g.�q:�P c�ѕB�p���B�z=�6�6;r��x5"BpB���⏚��>?55�Y���K�i�aL��CK��f�l��b3�|$��D/��g���  p.�U-��.���E��e0u%T�f#�y�����3���)�V���?%�xHۦةL��t �,Qէh��6p����}���i��@�O�01��>fn��r�vCI���lرs�!���t�[7�aJELє�p[��W��u��8[� �Vy�ի�ln�}�����L�^�2����+^��Tăx�R$�r��
/Ȍ�.���� �ɵ�A5NΘ��9�Q�����Z?�ż����+_�7Z�z�=��`'Ϫ�;�Y�%�K_�yV8Z��F���̳�G:؅Ӳ�聈,��G��φ�g�M�����ox\br+�U 9i*r�-�J{�Xt�_�#��F�Ю�e�kN��,�3�{
2?�4�gIp����]~I��&莑�IK �0p�;Bi�kP��=�[E������w�b��^�~��������VS�'�}�) �_�J�t`�"�[1�9rk7�В�P%[MZZR�T��4��yL���<�Fl����k�������va�鈥*��;т�~G~.��D��u�wK�l��R�b��8�a��������\[m |�֛>o���� `!��S�j;�K���i�<�m)��T �����.��g�ʡk
�zx"�`Z��ߗ>Je�+�0�r�H��)Ma�_��2/��#��c$y��^ݟ�zc�n��8��hKó�"�FN�8���o�$�/�, S*]̨H�l'}��GO�]4rh���<�M�����K�,ܥ�=���n9Db%59�4�F���F,s1����Z��#�L�����!f�<`ʷu�����tPcR�Jg���j,����DV���#�{�B'r��0�n+���%��Ⴒp��r8$Ɠ�ĩF\�cE�-����J���ګW�ty;7��3�:f�2I`�N_�]Wz�vH�p�	j$']���>@X�Ufy���3�C���$�B�	��'zjmI3��
}�a<c�q�;�[CܻC��ͣ��]eD���l��&oUR�=������W{�64��T�ڳU���/MЖ/q�rʁ��R2��0|�h@DD�g`�����F[{�����|t���ő�
4?i�b� ���?K�F�ik2�ُV���^�'�ـ�v��[e	Ω�����O������^ L���2�5⍱�^�O�Ea�*7Q��i���v2����H�I����>�!R��a��87��1��$!�gѸ
e�-*]���q"Z	�^�	ā�1kɁ��f�y��8pi��S�aZ����q���|�fRC�k��
��I�˜@NWD�l��Fq- ���af�}g�(�؝��á�U���S gk���J	`ߌ8l�N�����{1p�n���B���e7�h �]�����Ad7=�<V��)���Mpa�}�Y���E@ �	�,�@G��J=�S.�,�~����<��4U�J#a��o��_sF>V�4l�f�^�PW7��"�R���F3Ր�(Ȣ;�sk�ҌS��7`q|g3/���������T���#)�||��}hޓ���*��� �rw"��J|��et@��aM�p	+��U̚���e�gz؏����y�1Σ�&k�+n���WP��l������y�~�VtG\��⤱6�� ��˕���a�{)fzT�_�y�£-�]���6X�r�ܭ9Ie {r�jP@_�@%[�r�?��_½h����%�yE�;o�\��S�|�F�.k$o�qd:�$����~���µ��y>�A�o��(d��(��ئ���6�୼Hc޹[7�I+��rr!�.��ҋ�˱ϸ�S	�m�(���1%u�5�W���q��Z_[Т�Ze��Aw�jir���1g?���9�B5n�l�~�X`��?
er�q�wLME__l�*�7%�b�7��)J��bl������K(�t4���o�����vq�vqX��aa�:Z�)��%�LP��a@�]���	�����hB1jq�K�X?�+#;r�b���t�-�fQ����neP~���%���L�����6O���+�Z���M����4��,H�D�D�LJ��`��V�~u��!��o
vF����*0~3�5P*�]����f�o�x����,�UZ�>=ųO��F���~b꥜^¦GwNΞl�&�8��Cf���x/|�~v�n5�㎿h�`&���'��`�t�ί�i Mej,�^..)Q@YgW�V��]�w�о���ŏ,�!��&��L������,x��� �G��0�`��(�ab���=#��6���J}c�dL\'�2i�u�!��c�L�4���.�"��':cf�u�=��ϕ��o5���Rh�o{5�"��*\���d���?U����#{.�Z�%<�4���S���㚰�~;�L,�c'�U�����Hϊ�DC��T�O���K����U�7�UM��ޠ$J����M䊗AoV:h"��U "��)�C��
�=)�i�봖����,t��o/[`��#{����\V�")�ޡ��{Ǟ��`��������~%9�x߸ޫ�ˢ�l��K폡��MpH�q���Ucԝ��S�`�z�]���k�b���di�My���e�5����+��£	��w�asw��[LP
�K�6�~���F��b
?I��r}n������B6;��J9�bEf�������u�'DVy��ug��"miT��ׁ�zX<�)^֬! �X�
���,xyV��b1���*9�l�\Sm����)7���6{��a��X��E]��Yhy�kZ��f&��
�Vz�3����*# O�뜈��]S�|v�t@#�d�1ɧ�SL��GT��ޕGQ� ^}��p�P�T�tF��UJi*�9�>�W4��GYȵ���ä��߳��-�+���fq�}|;s�Bh0	
+ǰ~�\����5⒕G�{&`M�O�����@V�@� �J8aq�q>"wc�+�>f��������/-8�)�F�Zgv�O��X�BT�0'5t�~ڸY�"�'��d�/
JS�;I��a�z6�C�fW8F���w*��t�r�a�'!U�"��}��� �4�t����X'�~��k!��P���u�ݛ�n��w�~4]����H�<>� ���r�LEl�P�79tF��>���L�!�G�)
�*f�G������k��?x�QtF���T����0Zgp�!���Z�O*gG���)yD�=_�\�(�nϺ�&�'˞�=Q9�W`#�N�z���w���qF�ܡY�R�yٗ�A���Ox��W&����_��Z��@��I�'3e㬔)���N���)�PGƜ5���i|��EU�f�2ӶZ���sVm�O�lFZĹ|]����%D�͙i�XM�wI�D�	
����F�YqV2���3~7���^�����;�y<�F�ZF�k�7�����p�e�Ȃ���������F��0�5���$�}y�>z��k��c�P��%Gl�+�&㛄�e���x��Ҁ/��;�VX07Y?w�S?jfzb��$�*�)���
�|�M+��Q�xg�S�,�c����X����>Kk��nν^����t��1��р��  ߘ6�<��#H]y����^���o�o��f���Ǟ����)��W�F�2\aK����+yJ���>�P�GF�ރ��玲�an.=Y��2�z3�{t�Hj.�\�=� �N�M3ܡ=[ �>�� �B}���3���;�2/�)2}����.ħ�Ə��f>� 61��]���>�|0#�;����F���fB|Z��D
�a����7����͡�����0m�bSZ ���ޱV	S�d����I���&E6�VH�}U`�i4|�V��8۱?�����h)]��.�s�+�����o�/&��K��by�Y�T�>ώ��h�B����ȥ��K~z�ϣ��k��p��6�� �����PAzˮ�0��N*�ȁY�ӣNiG/�]���y��yX����e�Ǝ+	�f(�*{�Ί�;[VQK�:�����N/.*����G����$Q����;�����y�<�Y(�&"9^%d��C��C0'�-:;�f�ڬ�]��;U�E4A5���6����V�)�P�pvwٓ�YC#��p;VU��S������`3NO���~�sFl��F+���N�ڲ��*��E̜g3��6��彌C/%�� �	_���0К�8f;^���,���� �H�]�z�ݮ>�җ�s�=Q��!=�A�WC�brN��D'�9�Q��ֵU�wZzJ�>c��F�B�T?�����0�����2d^r���uV��b���� �1e�k�>���hPL��_өݔ��+�%ͣ_�t�r��dy~c�P��܊���=��WE�x�l�]7��h���>\Q����v�d�x�k�`Ul���l�ә�0�t�Aͅu�v��:L�R�^\"�;O�H<�/��~ܚm��l���o#�~LF��=��6��|��\US���]�f ���ol�埰-Ev��V�6&�3p���� ^�*�I��<i��~�0�Ӆ@�մ4�S���t�tY�FƆ	i�B9j�p�]�}�{�`3:-4�ҥ�w:��FR��jP�.���(�<�J\���
�˴��J4t��gM��>���ԗF6SN��'�s=j|��r�c��V��� y�#�~*�;h�$B���a"+�F�C�9��lE�$�Ai�ǣ��@�"1]�J&=�r���J���ս�������g5`W �&%q����ץd/�ũǹ/%pZ���pI���*C�~��Osď��^n@l/Fte��a*�pl��x��fG�S���	�>%�nZ���E���Ҁ^7\�ǖ�e���=-�~i���4��!R����6I�R/!=M�r�xl�W���#�S6�6��D(���������/f�S�.���1'b-�R��}���ޔ��긖�3��$ ��z�K�JU�K$�Z�Θ��7\ZR,�Ν��C?�^�sc��&ˊ�_ɲn�U�K�G<
�;�
U_]��Dd�hY�/��<����^�~��M+kd9�ն�*��i�ͭ-+�z�E���"��so��S�9^�b{Չ!�܁�p��{����i���Bݵ�X��,��3E�V��������?
)���d��*ٟ��?��p�{���=E�	2��'fL�$j��=�)3�����6q�xWV�������Xj�vW�*"��dig�J�ς�T��fj!��ҏ!�S8�7m�n��jXZl�g���k҈��� �9���x����#�v�Lio�������(iF,��Ѝ�v����}T[�$���E��d�>/�o�DZ{Y7Y��X�R�?ۙnQ�Î�f��x5rT��Q��rw%z�6ܫ�p�Đ͋45b������*�G�em���B�;�r�`:��}��!1 ��R.��o+�&���*ؼ9��N�M}�*®��Cs��9��кw�������{m ���~̠���_�c�rwJ�FW���/�PG�ZQ֡�%�I���8�2��d�c�� �fu��e걙���D��aS���D���M��
�E�u2+����-p(�g��:�Y�^�l��gf�쨀���(��n�8�H�G�g*�����x@x 4����wW&A���R'��!��z�h��2���������&�o�#��nػ��KB�V:$]R#��P�	��j�i��V�N�",�+�e��������D��F���4�Bc*¯o��4��Jj��6SZH�R�bی|�����S�W�A<L��d�L]dH}%�I}��(�YDb��f��	���N�0!	tj���s�j�$ohUe��"�ؓ]�;Ԅ��x�x�9�����h ���Oy��W"ֺ���9�ZeL7�ۼ�%-��o# !%Ȝ�3��xUV}�����v�Z�o��x�9`C��;N.���=+J�|9���O�M�N�&-�8�r����<��2Ճs�x��,�!d������O8ɔ9�<<�,��T��:��?)<����E�T��Ɗ�))Hۯ#���}x^a9grz�C;ߥb��1bN��8ɤ}%���T�V�F._�A[~"ѿ?l��'@�o �j�0�o
SkT$s�uͽ]9�f��X!l�P@ ����Q���J86���rE?b��o��� Ŗ�_�w�T_��*�I�Rcz�_���QK�B,�:��x�A�"MqG�X��6Դ�=�(�X lRV��2����dj�y��jf1�خׂE=8b��8D|{o��/6.`
�{֪��f/U��˳tӷS���2Y�r ������pr3��D':���*C����8����)�K�0�P�\��K��Qoy��,Bw�t��b��sNf���j�:��֥��,��$�2n!]`*lTҘ�o���}k��"��D�a������FK�
_Zn7�LQ�*x6tϱ�-,�=����1uP�3{�e:��P��|��^�@���J�5�ls����ώ�,�Zz��bT�1AlfR�x�����E5�ƹ�90Ѯ�EY�-;d�k��B�sPES)-.e�P��a,jolH�3��P�3�~�+u��1�['��oR}�D�N�z<-��#Ւ��h�P�7���"�z���J9m�R}8�Xn�/ h�����wo�ݫ�eZ���W`@��[E6���0B��C׌b��PQfV�Ѡ\�%X���Mq���:�M��,�[~�jOX�w����G������t@��:W��>���Z#�U�é�H���ec��lnp,u�S��M�q�'���a`Ϲ��=��o3ǂ�i;&z�Ý���V������d<a���5�S��"KA4��`M����D<H3e%̷��G-�oؒ]B�&Y?��:(�'�fP�T�G���.�����}1�&���rX�ٖ;� �o �*�� �)Z� �]�nsɧP��젏K=���7��ӿ�
��o���D
z�.{��s��+O^�כ����x���ȿ����ڱ��A�ojQ�WN#��Y�6Ü�+օ�s��
��,����`s.E���^E�"�0�(� ��V� [%x͕�Y{"'��9������<����r ��dt�c���0��g��[v�؀Yj,jZiI�ò2B�I�����9C��n+�S�d%��9YA'c��u8���ﺒL���WU���7����߸D@����0��XHP���:�7P~s=�G�OI10�Rj$�
����T٩p�M�w��ʙ\8�aւ�[�;���Z`KU��E���H�_��P�O(s�#���pD���J�ũ��k41�欸�:��i��Z���� ��,|�j��A��)H��&��"��`E(�]�����;M���B}E8j�cWY��������4�؃o��-`6�5�M���,�^*����㶈,2]����f��:�ٮ����,�^�~��/�H!.`���o��k�U���)���E�,����z�#�{/öW�(i)��BO7g�3����#&��3NKA��Z]U�w]5��\��X���q����*9\�OE�i����Lf�<���-�!�x�V8��L��^p�;��Zg�!���ٚ���\xs����aOǡ%��3��D�D<��mp��F=;WM�6�v.������5<2���s��V��傥�
K��v�D�`r����2g����:Ǘ�c�
�&G8�\D���}U��*#�S����{7�����v��0ѕ��Fa��P�,T�ܫai�{�̨Upu̎�we@b����C%f�7��b�P�����h���G�(�J#`NR���d���[�Ĭ�eJ���'�������o�bݗ�w�.kq�@�1_��S��uM�M��3�
8��O} {5��{�J!���xg�b!��1��NK3�X^ˢ�o�˳sǭ�I)������Ơ�N�����@<��;�Q]�n�_xa����І2���W>��E�M+��r� +��3�v0��S�
r�K�E�pF#Nry�^-���i�q�=%�����!����v�7��Χ�<6�$��2 v�u��@/��SXs\v��8T�W}�m��3�+hܯ�{�?���\�89B6L�A�8W`Ҽ�*�s��MfT�^��FMÆhVý����D�"0&���vf�=�tL���l��v;�ѓ�{`��ǁ��u�~��	�v���e(z������N�!a(�"8X�Öy��el�'�F+^��z�Y��Y/�Wj�M�b�NA�8����|sY�d�Bɱ��e{�`퐵i]챏x���]ͪ^�z��k��������d�{.2kQ�����M�@ӟJ��PkkCcR�5�y��(I� Ν�Y���8.�C1)�}ei}����I��'�nuK�{k��.������/r)����,;*5 ��Y�ݍf��*^k����
/���_
��m\�q0R��aX�ߋ���*�e��g<�B���S.a6�&G�Խ�Ɉ��bV�5�����4/�L�=�B�Q+�.�(�h+S���s�=�SP�:�CȨ�|X�Q�� ��<ml����~_�1�����k��$�1a���rlI�_���+'��l���/����ˣ2�8�˜�Ղ���wpox� d{A���+C7Z��U,AN.��,���\i�]$��M������7�/�f1&��Μ&3�W�|�zCL��w|�{w��3�e=.�VIj��X�hv�p�����3�).����WXs{n�\i:��av�JAM�Dk�j' 葡���`���J��<�<<=m�U�w�N��zL���H{BI�K�}n��˴��L'=o)��/�,����C&_�VŘ~����F	�mS�I<z���+��D����[L�iby|��,�D( �w��������L��h�n�SN����j�.�R�T�[C�b��^��4��mĿ|/8���\��ޘ�x�З�z��:z$1 VJ�����ni&[,@u�>�����/����?J){>�9�e�ҺE���m��a�ki6����D���j.wf����"Ku�����XU؁�t�o�f���kJj�>�Ք���K����g;���3�9��ù�{�@�f�,��b;�ٺL}�/Oda�sG��)����I���i���Qt��Ia�̓#�5ɽ�&�l����$�e}�V��?* �B)��etfGA�^p8�^i1��,���N���7ݦRs1�)3{[��[��F�#�����uAF�@���#8'K��Vae�}K.�0�e7�\��n*�2��8��U���2Ig+=�&�\:��ɉ2���8��]F8��Yc�~�ҥ���φ}v+]��ڨ���5������ ܋���?[���o�����n.�#.o1���%[kj��.L�$}ȼ���-�r,An�@]�mX^�Z��	���-��3u��
)=�cGe��
u�N���f�;�п�4s�vu��z���}ZB�i�b��/�<��p�Iv����qh�P���u���O�D�喝۶���g�G-v���h8���I�n�fE����V�`��JC�h�P��8j�N��^ɼS��f��ř���z�%'�������C��� #d�"5"��+k�+���p��1K��S�$�m��Hiv��q �v�]�������Ķa���-I	N_�fk��h�E&�KL�ǹ$[9�ρ9_�dg���I�~�c��X�����Br�\��ѥ}t�����~u��:�\��3Fd���~�U5�#c]�������rx���s/�p�P;`�35Q����e����{�&���*o;�a
=��OyvL��Q�n���{�^�fWj5�_��Y�u�;b���������ъ��9j�Zg�*5�[vd�K�j���7�֚��`@0�#G�\�^�^�����m����ۓ�2qz�����<1�L�W�D����[h>v�Uj�7��Kv7LA*K!�0;_W��Xt8��=��:gzQt�;<�0Oխ��,���L��	���A�~cӨs�GE�%��3���Fe�l�(��������ǲl��/EV�xh�u�{�zb�yT$+M�����Ѫ�N��Pn�)��$sƓ��O�vd�
N���4��D��j�F �&�(PW�5�/�(h�tb�Ӫ���d��8:ണ�@����i�F5{��L{�@"P��N	�ꀡ��Q���9N��H���m�s��$ D�z�H�n�GP%BX�&�d��1����!q��8��<�����\c��
l{� 0�W�{��;L=0�m�Z� +��	�#�${]d��L��.ʏ7�њ�~/e�O�R�]��̞��5\���wɖ���r�y���.�e�雓�� %dpU��a>3�k"�	`y�e��p��3�Rr��#�-oD�<>0��-���?�.��#y<��X�ݾe��J��`+�⯃y���W���G�L��-!3q%ں����z��bU��X�,��[��Z���:@�JlM/���c�j�8e�WS,���vik?�&V�Ŧcf��x�C-���"�9$q%s�6����z�H��IVK�v�p����E`ڛ3S����'�'@�+sWW���ڳ���)  2އۃ��S�57|x:}/�0㱽�w���9;%P.�W�{�����Yb�>{%�@�Y�z-�r"4���1R�؁2C1Ziy֛W��P��_y�K�5W0�\���5�����E�0R��G�S~���u���{�Ym�D�~��,Mz]Vĥ��U�RZ
�\"�7`.�j1�: �\��3�>���e_RUś`��؏[J#�wS������·�$��PV�)�I�<�@��d ����������%�Ly��>�5'�rc��z5��w�����������a��`Y����+������2摠B�#=�ZңN��G���
n�[�p�pLl�"3���GҪ�\�=�z{�*A2ذ�d�/���p��^�r8��(���``C Zm/�f��߻e�ջ^W!���~���\�����Ϳ�F��۵�y�}~k��7 �<��������n�^^��_�F�g"�"([���o������#:n�<9H�y�m5G��C[�~�\��u���v���i�Xj��'u~�O;���^��>㿇���*��e�$���,�z3�yZ�Z�����TXE	����U�M��'m��Ts�~"�ȕ��ϐu=P��㾓��2��h5n�)���u!%,�9���U%Ĕ"��ZqkX�;��*ؿ�p�)ͣ��N�D:2� l������T]�	����,��~aևP��j��6�Yp�d�ٹ?6�ǵ��\4.8*��M�7�������1�'[v�fEv+�J�]%�,8������7zy�6��#2Z��y<A.�y��������J�ϭ�����A�rW����H�恵r�|/*��u��OJ��ۻ����"�Vf��	��7�k_���i�ʛ� �ڸ1�T��h~��[������!_�<K����$�lڑg���f���.�|�#��R�O��w��v�^և�Y�T��ʍ�je�2��xB��	�-n{�������W�/� +�J�s%��5�}�Ӳ$ul�}8��Į�Q�{y5 ��&��|�l�6h/�"7{�ȈY�*��d.| \�,fHZ���Z�k�e�8�����}�F%Ky{����ݰW;���5˧�Oy��ɳΖU.����~o���*�l��E9�xyKV�ʾ՛������Ym�����p�B}8�I��E��έ2y�]!����@�������	"ĝ�I���Cg��E=[��iqa҂��uvE!����r��Q�4m����i�y�0E���(��^��&h��}C������ۮ8|�B��7y�:6޷������8�o�g^���k����H�7^X=�U������Ce�����u���{��̹e����\�-z����Ko?��{hԋ���7%����BW�-i"�6���u�����{�M�%;��C�8���NgD�N��3���]��vĹ���w1�a<��!!���j؇'�0�:"5�iF�����^C�s��j-q-�Zf�fP#��6�b�<��D6���=ev�I��Z�d�����d7+��C�m~���y<�{�\�}r:D˩,1EQ�2��Ӣ$�)	Y� ��e��)[����M+�-��ӡ�`��6	31�`0��\�"u�ݿ������q�?]�1���~?����,s��BXq��}a�7�W �U۩�rŪ=�V��8޵����8>����wy^�j�w�u�u��Ā��?��Q8�7�7�9�o�3�<ʉ4��!���4��K��>@³l
JkL��nj������K���G��5�J]i,��t�i���b;`�h����Qkq�פp�Z�	oK6�̈P��>+�{�ԩ�?81�XM\�$Oǧ���p�r���� ��$|Md�����_U~F�Gm-N�8t%Z����e㡟�1�x�^��/����nY��:����/~G"b�L<)��O�e�]�<= �2�)#m�F����X��]������oN��g��\oG���w��6����-���6̾ن!��G����V����&���Y��QF��w��	[��a�ؠ�W@��7��E��܁=o�*\9�$��F�_�8~s��%)��/-1�M���sY��=�����~�1� _����K���w�]��Nߥ�вu@ٜ#���]�	軔����\�F�P��B�s3q���|-����о_���� ��^�Cl�lї˅���|��^�\�u�Xq�=Q�M�D}�K�W ��V���K_A߅�%�lUЗ8ޞoկ�c����
U���k�+�o�Wʨ�;��)-,����Wo#կ�F�u��w���~�']�.O�:��b/؃�G5?������b4ӛ�eH���qGoWN��D)׬�ެl�V9[ן�e�Gy��/��hL�)�O��X�>ew]��������k��dII+}�A�ZpMJ������<1��>�q2��-�k<�	-|�w~0>>y��ҡk��5z�M���E�1vQ�f&�u�1�veD�> q?M���27��0���2_�z��UȡI�#��]���m*]v.h��@cl��WZ�4$�� �挴*���XVը~��w/y�{�?��>5�^�{Gb�Tm�����@/ѡ���h�����=��;<_�!Pnr�.����L����C���Fn����-�Ĵ�cy���w�:{еIs�E����![2B�$jNP�t���7h�O�?��"Ϧj|�}���z+���z�Nv���Aw2�G�r䘩8
�t2�rGSu�%��z�^�q���H�fq($%gt싍�]�o����Iy0/ډ'8�M�\�3�.�N�z}��јc��{�IiY����m���UZ;�d�Z�k��H�}�I�9���r����3��NF�2�C������]�a5U�!���� �n�Ӻ/��ເ�z�)ǻ%b��V�E��!��Ul����Wz�4���9��mNۀ����づ/�+�}s�4;�n$�Χ-��ؑ�J���ʡr,��o��ZN��=��n��s��_O�]�L;���Y��g�΅�$�,��M��zx�n��MjD���XSVRI�m�x�*Q��t�,����s�=;�c��sKzx���c�Oy���9ͱw+k�ʷ�Iq����o�>��G$8�vw[�S�dj���i�����\G߅׸F��c-V��a���ĔD��,��ͱ��w�Nj{�:�y�z*��j����y��o�N�ℭ@�c+�{��$���8S<bSMO�|Hݙi��}WAʢ�oB���:���]4�����D����~X��7��.��;)���;34�T{7���ɇ�?�����W���(�)�N5=#�2��1ʟ1����w��5�I�9�n[Ny|�]��X� !t6�!��JbYM�*B��%��n�}���ܽ/�d�I�S�m��U�8~�H��S�P��F��e�X0�잓����OZF��dOPl$�xݣ1^��+?�z1Wu����6H�Ϊe�ױ�.,*Z��K�v�|4���L�$I%Y�imj�\�!�>��[9��1�|�dIѡf�dʃ���a0)m���08�V�>�33��S3�ĕE<�5U��&,"�;�vX{DP�������InR�g��K�ٿW1���/�(��FF�d�ʚE��CO�e�_3#p*��tt2s����.!R+l��b�UP�_D}^��T�	�i�fk��Tg�Y~�|W)=\� >�%�o��~n��<��I��������B���%O���+��d�N2-��{Y�d
B��M�e���]���h�EUX8�2�$��7�W��+���w0�1je�W�{�#ۃ��[4�Fy��*�`ř��H%]�u��A�����^Ad�6N���^
Ew'U��f�:��$�h�E�z�!�Yb�ES�j�`N
��B<x�{8v�rC��j[���33=]ባ\��)�QC��v�/HR�T��Jm�ma�W��`�=����Blx�]�g�J�Cb���V`��-�D��xo�J�	93�[(��R%0�Wx��
5��2�E�'Do1�K���?��5 �ٙpy�u2��y��$3����v�A��7���B���V'� �> n�=�Zjb<�?ڗ{�/�>_cWAq�M?���:S׶9��t������"�S�D�N_��~R�,X�|fft�,	�/�݁�2)�|daoI�ߑ�1�� 5kx}�A��!�l�K�#�� �U��N�A������$�#s����?�z���m�yn�� �\���	���Ī��r:X+�/��"�j&F����y�ow�U�g�G?
G�Oa��8PKt���	ƙ�����^=�u���|�v%��n��mP��}���h�c�����.��v[;��#��>�=��*Q(g5�3j,J����ىK������n���s�2_~�a8a5�ϡ�o����Puy�̫���d�ۏ��T�-ܹ��G-�ǵ:��"K��]o�&�/8E��T��O�WW
��"�C��_���x�Z�%�,!�!޲�Qn�i���=��>fR>C�,�� ��P���(��ns��u��2�q�� <Yo��PTtl�`��q�E���	lgݲٔ��  {B��R.q�GF�E�������qLZ�J�ڡ�3�k��۱q��0�f�E�@�#����BH#NG"���E��:���")��	�ai"�N�.��T���� � ��G ��VY�7�Ќ�V"M�	1�ޟ�_�|�U�{v��P,=-ݖ�+[�0~���I��0v�N�+�_�>�I��+����Bܞ�ۤ���K�Լ�m���~���D��z�3d��&$��HplI�Y}3Ϯ�N�6�`^hH�,h��)s5�7�x�Ğ�=�f������^C"�o=�l�;��Q��:��s�" ��o.ȨQ�.�%���یh1R�n�Ffxn~,j����Mdz
����J��4e
P۠�,��7yi�^�ɑv{��iy&��n�"��{?9�&������㋗��:��c�.���ne-x�D�"�B�Ǻ�s�UB�P�r��A%�ᡃF�6��d��	����;�^�S{�����M��r^���53i���L�s�RH[����O�ׄ�O�q����2hĽ��MVE�ȣ҆v��+�/����~�k1���"8)�H����1K$~~���?���!�Zm�u`��_w���"�,�M87�5���a E�
�7��6Jp�`�g���|?Q:^��aE����r���C��i���0�*�3Ŭ�e��z0fv�a *��\-m76ڧM�:�)?���\쏁�4�Zv_��Gw��9w�ֆ@������w\ߴ7�ĝ`qձ�U���� �i��?��7��� ��%=�>�q�Ք��t��X�rX��&|��g������>/^�jcʮ{*9���Gv&�O��R}@Z�{�]�m�E�Z�=�X�y}jql�J��R�@���!�f	e��U�O}�����:�%��O�h� d��r3NŶL���̟Q� r4�^�:�uO��9hu,E�hK
���!����s�%`I���� �]I��f.�|���d\p����:[�o�s��Zo/��=.��Xձ� ��t��7�%{��N�S�)��]����$z�٥$cH�@Ћ�P��`���A��Sg�]��.�Ҙ�R2�RD��3S��Yn}ei��肟�C�9K�Jٳ��̫c%��a�{��n��ؐ�ϟ��c� ��7�oH�>��{�vq�-�_�����B�sQԎ
Y����n۹�!��k<�]2k�|ui����kqRچ��)�k�o�Eb8���4]��Ǭ	R�/�
4r�5�ه8��LT�AB����A��2�A��&�����(��G�)s������_�f�����L���͸��=P���ex�o���@hh�qv︺���mV�se딹@��t��b�v�x�u��1����I ����\�U �T!2vJ	� �b��$*�OޝPIC)��#�Y�FT2�$٣1����He��v��}���1~|�����n�#�D�Ő��E���#�۰
�u����C�v���j�.�{����g�@)��!*�[�|�kK���i�ӌO��'x(�L��N� 0����vnʒ��|��X���,�Wɜ��Z�L�Sk�	���s\���}�(��*R���iC	���s�oT�궪-s#YN�K�h�ެ���na��p�{�,��v%̾2����!�ç���ચ5�K�!j��C��-�Ý֮����C��l�VN�zTO��PE�^��Hʲ��U�a�+��v
(iB%"��?�FC�!�;�-��k��a�;�FSuf�#7��EG/_���A����Q'x���s`NU�L1��`�LZ�y�^V�w_���t���o�fT�
�m�Hgi��z �K�tJN��Fyfp�7
��%��v����`������Xu��]�܋�rz�(b�[�}JY�AZ��^� �z�����,�o�di�����ODl,�?f:�CTO��!0�� >f�u�/�A�̈�Ӡ�a?6���Ҿ����hE��	)�fͿ��[z2q�-��Ƥb1L-�hN��[�xh�E��J;� �y�mF�QU���..�/C��,�{�w����-o�|�"�8�
�hۚ��  ����AϵM�}�|��z.�t�2�sd.�!L����Y^X�$�Fo&*6l��]o����7������x�Oߕ��o�.���)"�'VR}/h8��)���Z������I��<�[��e��T`���c����?˞Q��7�i�o�M��p!8VM��/0�~j����R��QA�* h@GH�9�g���ʢ�W���^*��A���#�ۛ٠�[B��z����Yڇ�(��o�g �3�6.q}�is{�����TH{�v�A��B.e_�X[��F�u�v$WQ�-I��M��c���e���ԧ$�4�����l�RF	�:��?6��Z]kF}�<�lW��̵��NX�U���ow�B4��g�23gj%C���6��]�!��'�x�l�$�l�ոv�▶���W�~;�k�`gf��٩��A�A�������R�É�)3���R[Qs����}CȨ�b��v�3�Π����:3V�j��]�Av4*�f��1�\0�_`쒓7�~������$'!j�)���z�>�&O�đ���b�Z¹/t�Rs��>9��]�<���e]���o��
�h��<a����U1}��I�m��x��������ǃ�2����o��d���m��E��ֻ���s0
_C�J*�����^+Ց�uy����ټ�cW�e�M�kj�Kk���Hk�2�L�+��w���B6�z��(��>G~)`�~��t�z���UO�.�aH��_��P&_zO��:�|����:�$��6ysH �[R�Rv`D��W��G��_�����>1��Nk��?�Mi��DT�m�C���-y���3k���6l]"=���!qV[�KR/-��)��Y�)WZ7�ϩk�"�x�A��ȡ?�p3��̠E'F5PX���mz�~�4��O��AD{���_� �mʐ����:���a��E^����L��i�}�����v�9OI-nH�׋�k��W+�܁��f�=%���e��=%�qB����V���DK�F�@������)��ݬ���M�5܀��M��v�̃v�v����L��=�n`8��t���0�-:������h���ȵc}9�bM��L�+��O�TjUpő��,�}�$�/AU���4��B6����>H�c��\���W4�W�>��z�~�^�q8��n�?-�3eqs�߉S�#�!O|7<��>�T%h4ι���zCY�#��k��O;F��>>�-I����?�e�|�^� �;��������/�{['zD9,<�s
�}�Tr�ʡ4�Xo����b�$� �Cn+��'C5�������ќz���4v�F�k��J����Ʀ��0��z�t҄k��d����-P�~�G�c���,̇�¹��)�HA� ���a�7��m^j�
6�Lǳ,*���=r�b�C��	HVc\M!Gbf7¢" ��{����[Y�� }ZB����D=�훠)����(�d���x#3�5A�*�ˀ�N�Y�jrўO��q����%[bȁQV�o2��RU�ӂbTĭZ��:կRꛘ�Z=ɛ�ό)�Uu۷p?��Tig[ �aiW7o����n�d�P�p�If�Y�6x�}�
��3��A��}2�^-�?]2�6Li���}����SL:��-c^׾�9~S��gNr�&���I}�l��ô�)��(���踵�6Z�4�H��.j�nMt՝f9��J���$w2�h������<�������;$���fٴӓ"����f=?�hG�9j�.�%sWvׂYz>���	��l[�U����0��X9���~�EC$��� j�Hku���}}1��S��۬Z��d%�E^]���Jgңz���j�f�1,�=�b���dĔuoj�MN9��L�I|���	��WC�G�ҖeL�R�t;:P�ϱ�;�PX�d�j�����3�ֲ�{5�h�7GQ��,sm�g���ݷ�mB�}�4�l �Ͷ�<�Pu�� �]M��x���|i�D-����.�C��bs�����+SB�}!G(�W�$<�������h���`�3��U��~�u�a�����6��e{t�"��ꨊ�M<|��{~�??�'=|\��VY��P�(z� a��q<0^(�"�~sA�I��p��L}����?����,�H2v�2H��]��z�u�����L��OAf��H{w�,{\��E�����E�B���ق�\�	�q3�a6-�M�o=<��!����p�	���^�<�z��@����1��hdy'�1+�ar�X�	u�zO���̬���j��!���a���s��:�V��i{һ�PR�R;MD��	��M��L��:K�M�[�&(���8�f��}����,���a;��x_;��_�&&C+�'H{�4�j�N��,FZ2Yyjf���/��p�dI�u�����^��]H*`�x��:�Ȗ��_b�e{^+>����F��O�n���ݤ�������"H7������c��s�Mhi��e}��b���RCD<�0kyo��a��PD�����s���g�}� ������ْ�b��~ ��|�I��p�8�KZ_��ۡt C�i_'�G�P!�A����>p[,24�z*u�$��ޓ�꫟��ڹ�c�]HY��%_�T�6�e���/da����qܑ�V�e�i�;�:Y<�5���΂� ���-`�=�������M�gi�����qx�5���W��Y�ϔz�;?<����㲎8]�!$�_��af+8a�T�%��1�A����=���
b4����~�<�q��Enz@���H�&^I�s!�z�^)��ؠ���,.4p���f�[G��X`q��~�@|۩q��jkykv"O�\)��{�u�Ȯ��|r��rz��@z��i�G�&��-���;)<��p�{���UZ��IFQa����\��忌1�a�y)��7� �=���\�˶�d��Ƨ���]- �?x�}ȹӻ\oHX\���+��\Wt���%?�1����2�%a����͖l5y���b��ׅ6�X6k�%5���ʺh�nY��Y���8/�lr9¨я�8���o�3�P�� �sY���fI��8	�	+N�}��
���?�v���`o��Dk)� ,�ik6��?˸����
�ٕ03��lo�)/��B��ĭL�hO�|���)��Qk4?�Z��=I��Z�����Vʒ�� w��j���~zCƉ��R��lX���%J���ؒ�5>�ަ���|�I��z�؛�2P������sa�C������o=.��mы�� �O���&�鄾��=<���o���� (w�.V'��\:9յ�2"�l�	&�\�.8�7��1��%���$������q��΄��}?�	�ϿmmU8\s�xgVٟ�5���':-�Z=���})OA؁��DvK�6�=w�����J=H�PL�T�3���Щ�SOw�,!�9�%Im����]��[�q՞7�2�Q�0�k�xS�t��)z�)�v�bKHR�"0���7��[9E��#�v,թ�?r�P;h��bz��F�hߜmS�4��¦��ܺoRWp�_���г.G {mP���u��6��J�-����z����1���%fF��+wZ���c�]}�v�Tz�M���R�����b:�*B�m]�s��D:~5���kw	�mփ�ɑ���"�5' �8�*�#� ���ayB��>�&�>�47Y��y�n|��9�,
��*���!)z��2�4FrjX6_M0���C�#�`��d�Ӎ��<��e0��#?�:��.�?,(�X��N^�t�QhYM\*���p�x$Yl�c>�u�4ְ�z
(T쿨5�c	=��W�2̔��x;�����!{SYo�Gfщ�[��P6���|�rU�i�N��z�6�����h��I�]�%&m��������y�P��Y����0�Z Kc����|x�_"�VU��R��f�|��������}\Q�O�\�qY���L�1�v�
m>�)	��h�2�JٰJ��Lu����!�M][L��.��t�LhU8��=İz��ͫ �e;I �l�ԶX°F f�����l��Az�6��8u���A�0ZF��u�Ww,�����Q�$l��~5�_��rPQ;�Xq�x�,�1��%��~F�C�0���!,�Z������ʑL֮��n�P�m�m�̩�k� dPܗ]�ko��Ӂ� �Q Z�j'���UDs��ŧ@�>.��Iv �+��lMy:�����4
�Φ���D���}�ч��+�5�*B^�+^5�HDy�rF�陋�/���Vh�.>=F�W��Z�ُ9�g��]w0WM;�i�M���_`��F�S/@<&/���$�`��vk�.�{�Xh�߾%�L����\�Th�آ��xu(jK�Ȳ����r������R�����I����Ч]�����h5������~�� 	ht��װ[��$r@�XES���b�y#�QmП;Me���#t���Y�g�b��8!	�[��M-S5֮�n.I�P^W;�<46������Z�gJ��G��̓U�dwS��RROW�컺R`
+N+�i�%A57�t�k��"��ϸ� �������xu�^���eC��n, �1I����י�Hrq��2/J�A�W�����@�y�WѩQ�{}(�o;/���;Bˑ�٬ѳ�?,�u��g!8~}�7I� x��s@w��W�%�����܊��.dU�Y@��T�ߦ/��ި�)�v(�jl%�+�
A+-��~Z� no��Q�vq�i�v(4}�d�㫯�ұ��xX�b/�FA��}wP2$~�"ĕ���x5�^��yg ����dNڀ#�jUG��pcB����K`����6(!��C e��:�<n��\�6t�M��V:>��)���Y��k�榺;d
�~z��'-����;���Z��O��A��S�T�D�&��F�X�Ҳ���֧-��
���d�����**�|u/��o	����zT��7�RQ���j�ײz}�o�y�>Х�˶��� r�&!�ɬ]Y��	�6[w�� ��?iN��ڊ���z��ͺD�� ���#G}�͗�UG����y�[��E�y�/���sߪH����2��1�l���V���Ȟ?M�<��VhNC�̝1�;������PC�US%��S�i�j��w3����� ��( ���[��J\���OFO0�3��c���`��Y/�������AC��B����S0��]�(��7KNULڿ�>�U�l?-�{nZ�g%zv;XM�����]�����(����*���o�@ƀ����?��d9/��o]�~W��LEk]��(�%�Λj�'5ib�IiO����Pg�f�h˧ddY븝ˉ�i[�Q������q����G���Fz��16���߁��
�K��Ȯk�w�9U/~w@�XXJI�Oux8��g���� �eVg��4�$pvHA�?/�����i�����4���0W@���Zj{}Vj�V����sq������уW|)�`O �l�.to����dZ^�����[W�N�pe����?{R�n�>%N�$3"�J���Ҵ�)��c��A�#&%ZbjGU�H/k���U�x�Lg9L)=|��O�E(�i����V��t��%$oV&q���P���3�0��в�m��%bY�}e,8���.��S~.�%Y,T������Ao�K�&L�C�9L�ݣd���S�|TK�%�޸�9<���7M�8f�è4Ԁ�}�;���oyX���zCL �3�~�j�]#C�;Sm�H���:|DuCI@*�^�7�m78�m�����r.���+VH��� t��-�˦����>�,��gi����g��A	E}�qj���ҩpcl"�N#�Ks���s(0���P�dm��w3����f�`�t������/,5�f��o�2;��ʘ}��FI,�(oV�d$̈MeW�*�<C�Wˠ'%*P���_����u��Zb���g�
�L�t���?�P� ���WL����m���{c�]%��-n���5]�/�(nOѨf����d�oO�?#���,Ma�cque}E���a`��픣4W�ϲػ�C;y+�]z��<���z���94�p x�b �Mc9��~>uH�-D/����|hyv�l��f /� �5�^<Λّǿ�����F����x8�Z*|�E�!���"j2;���s����������~�ku������lHN.��0�{���4����)Y��C�!����9Ⱥ �`#t�/B�"��U3O,��]�ɰ�x!� vGkʕ���އ�שHǔo@Ke�ga���a'~*��Ě������7�#؇��'u/��W�:2�=������ă_<u(��c�>��'ypf�"$o������i���`!�_�{8ۚ�ԗ�v��dE�
�Y�@m+u�m����ͼi�����nm":d�Uz?s�e���Թt0�ҘD)�F�u3�#�4���[���\,�c�u�X�H��P*��`�����WƄ�w�6��n��,�7aY����tf�)}@xt���e
~_<�n�>u����{�~��BnyY=F[�f�[�=1OQёl49Qr�q����G�0J��Q�}�~z��`_{!/�ă*����47 u@�g��֠��؈�D�S��BcV���@W���剟 �}=��U�{�*�,A�V;�ց������+���O�]t�F�pFL�d:� �5uc w��&$�< ]Y/A�H@t�[
\}��B������h�~�=�1H=��Q/���V6���9�6Զ#�D5���z�ű�:VZw�R�Z������s1��.z"7UWa��F��)Cn���E���ϔ�Hp�j ���q:b���E~�?an��������8�LGB/M񧏺��ܦ��M�����ol�O.��cRR#����گ���)̤�,�tS1���W�u6��� ��]��&R�z���_�~�����)���)w�.����̴c�*j4V�g
�� �����f��Om�6g��E�,;�O�Z���� X��[^��7R���. �*�t_�c�#9Z���ԧ0p���+6���)��N�H�s ���c!A�O���~jM�BDά��r�	x���Qv�U�뭰�U���ڨ�A2�㫮lo�P�s7�g�Th����Xj|���Mh# -�"�?'��󍪾v�v�}k
~��~�懶�^F|���xYz2XC�!��o��u4�� ��o��u��u��|p���\�f���Z�~z|$����{�?�?p��"6k>X�����?>�ӺK���a����p?�~h�?\+>"�P�R�K�.U�y}���_����V�D����������,��h?J~E~(��s��շ��\+*��z��֏�$�L6>P1U�}��K}Z����w�
^�lJ_�����S�K2� ��e����Ty���|킩�L�9f��q�a�vi#z��*4�Q�����i���e���5��C?�-`�$��gL����A���w���q��p��Nl�P8#���;n����B	~wX�Pfm)�G<���6�Lx�E0���D�-��)��j�b/���UZY͞:/�������6^�XFCAz��&�Om��ε����D�aY�2����K΂�c^��=�I��{���K>�v��-.l\V@�bS��-��@���I���/m�?�.w
	 ��)�J�������$���8�/'�hsʪ���Vk�ƮCW]5��� ���ھx����X�-궉���}�K
�g�RSkܯ�M�$�5�r��Aa��1Z��/�
,�w� ���K��5�����_5�����9o&��LK=�g_�i��X�ᒶ��ӇQ�D�Mx��ޜ��-�^Ѯ�{�[��:�+c�U|�l�?]��?Up9Gm�����y�i�)�0N*���e6�cX�}G��7dF0�%�g-��ñ�vh	���>�\�׿������lv𻜖�!v~�*�S���\8$�T�0�����ս�Sm[E#sE:��N��&���u���m��{*I^o�ק��V�]|�tĞ�����5�7.�
��
DP�sG��R(&�<L�}p��&:�4���Dܮees��ݳ�"!���D�-������DR�{{��} �E'��R`�r^YT���V�l�Y`4�܅��a
?D�ȡ����l}O��)�����U�`�Mw����^_��B#l+4��u#Df�F����(��6�	v������\ԇ���p ����i�m7��sxXqʹ��{Dw����j�/�^�<L��j)e���Z��^i[�w ��uF����X��|��kZ>�.� ��i�Zx�߶A�} �� ��D���[I���xZ��u�V,V���@JI�^����=�y���O��� ;j�J��YS.:�->���@U,V�w���5g_C��Co��Q��4�װ��$߬Į�ٌ�G����b�،���6L7I;pD�Ξ�Se���/�z�`�l�l)�&қCmO2Ej ����l ���rњ����2߫q��/A��f�b�U^�a�>���|���z>�7�qr�TLm7�N]҄�@/�y�2\E?�'���I��v׷A+�$�M`�������*��]����@}l���/����l�j*��8N���b��^���0�p)k�sY
��ο�{����Y��zq���_�|q�h�Z��ϰ	}��l�?߳'��;��_�_�-�u�]ge�|����8[s�/� �3<b��s���PK   7��X�ة� � /   images/3c114b42-368a-4c2c-bdc1-509aa8451bd5.png4Zct]]�Mnl'76۶��F�ƶm�qc�qc�N�_�o���>?�^{,̵�<gG*+J!������!�H��~�a``���_OF �̯�EUJ�f���LF\D����/�������zje ��} �,"
^K�v6:
6�q3:* �6�@|P��FED8a�K�AM鵷y
6�9�k�q˓��s4.�����{b�7�sR�������r�xm����	5���x=�$	VI��\Ҳ��L��6E����ZܘTIy�c��4n����bO�������'z�<�Q�w�ڹ�[�@��p���UܧJd��ʑ�T&���Ϝ�F�\�|��Q�Ώ�o��������M���NIg~�5-K�??�-����;��C�Y ʥ�W�8����xڋ��G�K)��Sq�U:	RBt�O���eP.��rΧ��3��nN�~�]�%���L����9g9~�@�a��z�Z,�'���[��"@�aW(5!��X���d����z�-3�c6�,��T������P+�);�0Bg��|a1�_`�@~���b����'�D<M��V 9����-��\��:�	Јh
Y�P�}��d��ƭ�;n�+[�Y�{��9�y8���Z�������^��lG�k�I���o�]W[N!p�]/�Ur>���I���,	� ��9v��/�^;)F� 1���u3�UT�_���#����������ڟ\��ܫ�8����͑�v�����{Mw�	�ם�㳹�qu�c�)`e��/6:Q���/zɮ���� L�p�<���,ב��v���G���ڹ!��G�'q����Z%Y��1�]��ޕ�r?�)��t-&��]�5���� r@��h�y)v�;�?r`�D46��U?�F��?"��hʧɲ�gl����bŲ������O� _� �ƣ�n�1�5��T�<���u����d�Bm��JGq5tj��Xl>�}3s ���ےB��<5O�e���HS�y?�>�-nw�n�2�S��~R�q���k��k�$	UT���n|�{;��5;�y��Ñg�
����,r�vc�ߠ�Cvχ��1�����ٸ=@Iĝ��Pb�.&a	ݫ�&���|��|�����6���P ��i����u04R��pM;��.*d"�T���b[�4Be�\`�G>���z��̓�����y~�:�h�Ϋ̅*�-��􄒈�S�u�Ɛ Ih[T�U%�w�+�'{~5p�?|��wv��Y��*�y�8���5�p�j�k��&x�i1�I'!"�C#��Q+M}�/�
Լ��js����a#3�]�+*i�4c%���
dLɱ�ط���[��Ϲ�QQ�z	��+w?�w�xyt-�if��ǆ�	�&CM2�Y�D�Z@�:�k+Z�F`�=�Y��Ώ��]�,�ޘj:,T.DVy���7���!AE=��u�D�&;���A������c����H�6L�T����f������}&�5:|��5��FF.����7z"c#�Q�vvfQ�}����W�g�"��q+�ϲ���[c������$.#��x��ސ���S6�jA�Qx	�@�rG"��R��{���S�U���x`���x���[�R��N�Qw�\�5Z�L�h>4
���/�%�x�7V�u� �,˝SFe���Å��� ���v���!|�-.�oE���?9]Պse� �\��찾�db�`̢|�M�A$�s�?O�	�gw���%�y��u�ʵ�s�ړ�1G/�f��?�q߮�#�OР����2�حg3V�!��`ȳ����tr*I+Hǰ��s�M��̮K�;8;f��:��u?��j^�q�F���'N-".���Z�o�`]|���s�Ƀ�F҄a�I�67��6d*�0
���r���5zT1�c&��~�B!O����L�`9h�SV�9'�T�<~��R��TEEERο)%ï�,
�������j�����j6���z�-lgK"�ڢ�"��n0��MV*�e�~/��yX\&����[���f��fQLLLL�Mr� mM� M��U�|����#O��8���~�E���{,ZbF�v���J�a��h9��6� )���v�X�b��w�!L�u?���Jn>]"��;���2���b�N�"����\#��w�:�M��?S��?�ɿl5��|�����.����cL��?b���D�E������E<�:��r{���,��H���50��^�XMC�����d�	�_#�����A���6a8r�Q��o�;ڒ�������l�ۆZ֖:p5^ȯ�\����Q8�az�0�+�c{m4��[æg�|W��JYx�M_�.�j����s .�h5XK{��&��!�A��l�{P�Q�'@D���ڟ�y��ّ��|������q��n�d���c���#����i��0�9ԅM��n�-NI:�d$I���ta��̽���$6�<F����@Ny&�=�D���f�������z\��'@�&�Bl�c�RC)�h�����;t4T��]�1 ��6�4 
���P%&5:�L�%x�٩}�UUltD�+]�&�9�7��	I��e���*g��kb�4�'�=N-_1�/�Iqt���)��B�7/[�T�/���N�����ҭ����or�u;�Hs��p1	���&��t[k���F���G?�K���Mi;u(2[<�zg�T+c���*�4�z���J���*TԶ_��Y���^��=��D��1@����NMK
V���]S���,u&��qÅ�^�4��m?M�5�չ����&�|��O�>@�r�����72��]k��y�#�����+�W���&.�O�����,C�8o�D��Y*A�ê>t�Y8G��^�B���N�Iؿ+pq*���Dw���2��aH�hhp��9�ξQE�����>�|B��>����>���[�ya�����;84�lM����$����J%}��$-
+Ga!_��@wI^��IVlF�$"W8�Q$�I�}��pJw�M!��?�YU]a�/������W_8��苙���ҰP�N�6/z�he�������(�*�%�"Nv��R�����@�&��݄��Q�Y}��.ܗIʌ0��}�����W�x����#o���X0-�>����F�~��;�8"P<KV�)�"I4E7	�
��+4�r �M���TBr5�g͎���U����Q�Y&�g�-�:�3�9���K�^�4,p"��*6�J2[�0��e""-�!&^�\��6�� �eb��r�Y@�\��l��C���}a5"�Z�ʎaE@�KL��M �������F�t2�:�pA{����pRI0�$�h$�Y �Kd�K쥮�������DI��AQN�T�v���ɜ�R��׀H�M��/�PW�זv��D�]�Ѱ��,�+���I��T��u�):��de=�h�H��}�(���qK�h�!���w)��Io�C����s#���q+l���$	�~@�0�r�nt��{O��6�S�L�^���"��<�Vj�����F���<|�^ry��p����|��P�0;�1��*6�]��Nl`���Ѐ2ҝ���L��'.��B���oo0�dk��l���+p��m��d|	�ߢ���n��-/����=����?���W�����O���!cn��1��~�nڰ[M�@ 6�<\l��U�~�ol�D-��cZ-?e(ANaŒ8G���w^nmK,?֨����z^/��V����.`���VZmǦ�Ă�k-�d��g"�uڄ�������jLH���� �<�|^W�~R���V|�H��+��)�8,L߫v����t�*�o90h���M�G�/nޣX�7�;'��n�{D�n���F����9�A���ōy�n剌������o��]���3�O]+S׺�U5����}��G���2·�n�н6�`F�o��4m6K�l�
U��	��!~����%C��L�@I0��ﴸ@�-4���l�WO�b�����>#�p1	l�7�T�aH߆Au��}0�	W�-���N��%SB]l��6].g�}o��j�+���5-�s���^,��,�"K��{ c,�Nb��[�y���+4��~���h��Ԋv���#[��D����21$�n����8c�5�Q�ѥ������Ui�U��]�����g��3�` ��bEt�u��I����鶱����j��r�뽲��l�]|ɸ�8��4&]�s��:����_���/�yT�;��x9��!�0ZK��b���/�'�pEma�܁�E���y��Q���4)�����'��`�S<!_K�r�iz��G#��d�j[�������XG�p��l��e��|-�.�a�>��4�Ð�vޝ��_�o�������f�z۲�	��@���J��Zˏ�ƛ-�S}����\O�)�^��ndM�&��&믺��� ���.`�nz2t=�+�E��e��n��[{=.���5�wd�3�K�������»�4H�ۮ�X���1�:5t. �Ǡ�ş�m5Lgԟ1��`Iк�����p>���x� ����G�����^���d3��zI� �)���x��*g(Ģ�� ��"��&k������􆾶2u;et_r���8�D{7Ϸtl|(6���0CU��$�X��qfj��B,Ds���{<�I|a���\(&���4�=�j&�֗^6b����v3��u=�o���#���]d�1�������e8�Fa _���/I�wO��8�S�ߺ��?�_�Ϫ�l��Y�à@�_�m�K?�y8��yd�}��`ID���*�ϗg����n���B�jΙ�bD�����Z��R���)�k�*4 ʹ�>Ë� �$�S�4���tCL�5���y�S���ƺʌ/ �db���j��u[:�#��{���������s�q�[��b����R�3���܍����" �	��{)8�bp����
nr���������l*�*�h��`�;~�nX��o�f*�����AI��Q����.�i9?���oK��7�O
�Lh$���/;��q������:���>����zpF8��=�xC��{���uu0p6�|JIIa]�S��9S��X����r����,�H�Eҭ��0���Y�=� ���`���B��82�����7��	�|n���{kT<�N��3��l�PŻc��'��p�Dd�7%P�,G��~o�/����7�t��C$��:i�K�;<��
s����cw��26�h�ӵ�ï^e�l�Q��)����xG%����^
׫+9��A����8X>РA��7��R��8�������1��䴖���B�7k�]�Ͷ�-Xc��V�`W����/\r���z.{�_jGC|1^0��y�����9�eD��${!�Kat?���׹PB��0Vz�����t3���LB�s6R����;���o�?$��[��T�h�������E�ea���L�����p�\*.ǉ#�a��VM*�34@d���
GE3�H�&�mk�G�sL1�M}���8��"��G@0������C�Rʋ�n�_轤���~x�s�a1^gꭾ�^9���f�U̅���K���D�L�ewI9�k�;�e.�~���9^��#t�]��0ŷ^�
��������K�/L�455m��K���2��ٽ�����>�"i�<��nd�A�r�p���YXƕ��z�N���:���TR������V�o�H��|����D!<��Т �p�}�	����M�4�^����V�>�ߟnl�����w���+��5	�FD<֫���ȗZ�˵2�/������7�,ty����������� �ǐ4�d������Xu��ٖcBFΦ4�p��W�d=�+��={�����R_a���[g,���L��Mжo��(�6&�#JƼ]����i���b���_��-������@a�"��r$՛�Q}Ѱ������V��/>"dڶ6V����f��d��`csZY�ŶrA��5����yt����&�!��c�N|*�)#E�~6Q-�2DI���ݛ��j5b܂��H�.��q�1gLR���0�;/���ɀL���"�?,c�W�|� j��b�%o���W<��?�:.q��=n�~�� c*�r�D�q,�_�u�V8UֿX!*�؄;�7������U!��l:r[`�V�C�l�o�)\�K)��0�v�wi�y��	�Yv�]�}y���i@��d*:�ʐI͕.sb�#�h���%X�B՘�O�Ӝ��:�����G�)�|1,'�U�8�����N��:Z�$�����*N�A�i�C���*�gZb���C���@4���

�}f"��<��]��{���ֵF_AC=�H��ߚ�*z��(���[m�m�C���������9��d|��}��v��`bη]�L8j�s?��uy������ר��Ld�3�X���|N}���ÝLw�������p��siA@4��{�g�H��M׵�,l.�N��Ơ��[�7]��=)Sʯ��D�]�J5z=#E���b9��r����<%fZ)dF`��d�Z�C{��{�m/�p7�H)y��N �uW:��1֞@)�٥��z�"�����7��\�_�3l��w��"t��dG��ZK|(R�N��%%!9r%PA����-��������6�к��h���E����]UV�o>2Af,��p���."#`h����l���"�y��@S��*j��<��e�)�8��&Ȕ/R�{���jCmOG����?
�II{_ܜk&(�k*������`jh�iXG���l,��M�w�$�O���o��ttx��u>'8�M�����~�/��[y�6��v�E���&��t�f�����9F/����Z��{kD�~�f�JJ%��!��f	��=U���q����Xr@=���+�9��\�U�Lq�٨/h�+�G�~S��%��$�����.~U���X��,�)Q��$��UV��5��[f���쮐�-Z)�d�I���P��M���r;s���lv:��F��9,V�j�ֻ��]�������{Nl�D7e��{=_�F�y�3Z��޺�2Ԯ��X�9%�xT�մ9��tj��vE�$��~�wBq�\,6�5x�a8+bw��y�*�_��<M�� �X,'s$���;N=$�A`�W!鯁md� W}k!�g���ʑ�U�
�eC5+.R�8����T�'��ð��5��}h~V[x&`�:�i��>��e	x?���~챹��3r�O�"i2���`d'ʈ�^^��������a�1���f�[������n�OV�lۇ�0$|�p���T��/<'͑�2�w���Onfi���[w�سJZcG^
�#��>^B��z��'^K5����לG�RB���;#��21���/I���j��F
�y��|_�������s'�k�{�6 �Q��Y(�H(`����,LZ��4��J�1��?����s�^Y�+=��G���D��m�у�Q�Z`N:�R�5[��	zaT��+T�2G�S�� X�E�#�8���Y*�J�ac�
����8���G�a|����y~��K���T%h�#Ho{�ER�|�w��bL/��������9��h�(f��%� ��	��9Ŗ?�������6�?��-s�L2�E��f�	>�r��1�p��A�� ���	�j��ʼ�Ȼd��p�>��\��ǈ^�\}e�A���g/��/��~~���f���]a�=�-���	�1�87�x��p�a�E��~F4q� ����+C��_���#/�3qD�ԁH^��L�C��s��>���.{O�}�[9mJ�/��f�z'��떬�.aR�eh�AOD��by��αyp��(��
�S���u����_���'�2]\����l�*�>o���{�B&�z�b�ΜeBn�{�l�o����+���#~N�р�9�7�Oq��#�cLK��`Ez�U
H���'�"y�JcddtT��{�4t����0���Ip�"��O�_�'S)Z	�=uf1D��.�+���)�r����
	w�G*����*g�T�tw��x\T�rG	�Q(6�$�m�
�|zeT�����C!����`_�0��pN$��"�@>O�>��T��屼���T̘e�~���&����袂횰�Swn� �����K{y�n�%tlK�U��n8�����u�^�<>�-0{�!�!Nn��+�{m�g�S&U���k'|�����m�!��\1:g�LC�I�����5��
O�X�w4�F7�Z�]�C�|�[�� >jp	��,�Ң��Dh>ѿy|�@�k_:�F�Oy/�^?����8]��><C�oA=?nQ�����}	j"4������z��>7�
�ys�Q�+�I{w�������n~��z�3�}�L���M!t��h.1�?��������ƿ�n�������]�p��X���W�H=����u��2U��<��u�3L��ks4V0���+���Ԛ�'��f����۴T���h<��[e�}�������p����Ȥ��6>W��C^��ԑ�^�`�p�Ç��c�,"�U����ް�С}�XчըT��B�s�;`������=�c��ӧ��zi'�0"h9f�;��{�L�6]�U�����}Œ����?������F�<���Q(�F_ߎ �
�o(�<��-�>[aXV=�34�p���BFͣ!��Rs�\o����Z��z��zR�q3�}˿[;�[��)�����k0�M�l҇A�����{����t�o��g�jH�����N�m�[xN\��f�-�_�w�]��A�WN*u���L�e��Ó�r"O�9�[K��y?�k�FjK!�g�ѿ}��-5Ԧ�_�p@�����ݭ�t}���!3�ϼvk��B�8��F������Gb����U�a���w�����رR��},��'8�{��P5#�ft���5�:9¾��x� ��x��P�\q�����"Z6��F�;�R��n���{0�57�$�Ӟr�+��4Ň�y��`�d4��� �D�4�L"jz�H\dus�߼�P�<
�c����D�6�=����<t�D�a��L*���x�2W_����J}u�Ο	kab����4b�R�{�����z�!���`�}�K���ߜ+�3qR��UmE����H�EZ@OӞOe󀽚�R�e{�0"2�ze��*�K"4�j��x��|����,��5x�8C��"�����Qnu�]���h&6�U��m�
<^�vn�U��6�Q5��������	�f����	}al#��QM����f����M�)-�&j�B<�P�=�,���G;{#��:�HO�;��"ϯ�=���Ѡ:����Cϙ��ُFaI�)��t��Ym�qj~<���{�ӽ��y3���B�p�mk�G%z.5����!=$$,b�-d��e�����,�G�?=����I*�*`�*�*����J� mUs�.�@��x.���63;7$
z��*^�)��65��Nl:�j��a��m��rPJ;�svɆ@�9��U#�C��X���ڢ�m�������zG�+(���G� :4zM/Z�q[�i�W(ɡ"�ߙa�B����g6ח���C���H���b,��X���$�:��~�`���)[0���}�IA�H�{�d�27�VyybYp�°�_K#G��9	X�4�n�b��vgj=�EAMy#![�~�ZV��HJ%	H�"���.FMHv��;=e'Nő@o�x4�"JI��Y[E����Rp�z�E��(���J���]��H��T�l��NC�ҊZ�}��o�U��t�j`�k���s/��1Nd{O"��弧�J�y���޾�>*�W0�n��Y[re:8J�i���Kۻ1nI�׫�v�S]��uR��Іղ������[[/��OEU��ʰ[�FƧ"�D��P���*s�D[��B�l���}	g8��&E��� F߬�S���} �9�U¤F�����d��"D6:.���	0]�<|q�NZW�8�:���@�Ӑ �>kҶ�I�!s�o�8�^E�}��T��V��N>D����l��%�%��\�SP�(��y"P����u��d �g�+��o��(��|��A��WV�ڰ᷃�H�#1�q�$*/�"&��߾��d�>� ex�w�+jm�V������h�s���S��Cb��"��aA�v�,�ʒ�&�Q�f�K�Z���r���eW,{[,�&� �L��tkts���u2�H�l��'a^"���O�e$bh�y��z����#�r���%v�����J�sLFC� �+�|��98(?H���u�\B.�����N���+1I��_��&��A�6R�K�ʨ}`i����d���N�"D�uL�2��023�Z�a�h���=�B�iF��������� �fy����l>�ro7����h�:O��}{���>�q,v'��F�t��p�������,Y:�!c��Yga�tM�~6Y{ڌdF��j?�������z`֒�s�n`�5j.G�"�G���@>�Ó��KF:�J��u�f4���ϡ�F�>�]�v���Š�8�#� u���\��჉��q_r,bD&�v&7��.6�� B���.�e�N���g�'�<� �;O��%�qL��⟞t�-9��=�+X�n��pI�'��"1+�!��RS �oy�	�k�ޝ�ߝFs)�f
x;eo�QWw��Bq����C�!��^d|��b�*6�T���]◦T�KG�\`A�_�d[������,*�ތ)��-̒f��n�n��$�L#T�,�H{CK�O�- �P5�iE`�ᬾ
�TP��O�������n���G�(��
qIǱ��H�wC��_�;ϐE�4		�;[�9�˝'���+[��x����Xf�D���y�5�Tc�GrX��a�d�ϑ1>�z8����#�rH����М=|�̦ˇ_���� ��9Jħټ~?�Ġq��3D�-�өfbp�}�A���:P��i�=�v��\	~\�����p7���b$:��d�[箷 �%ʐ�ܮ��3]0�K����H�ĕ}{��Ps�P�Kn��2?df1�3����шT��
Z��w|3L!�X u�7���x��e�EN��T��9�Ŵ����AH:		�Ce�F{�������;�<�A��J�v�Y�\���n�|�+�׺�}	�.!�̇ëἳ��.E0��$A���'�_Pa�2ܭg��?>�
�й�i�ڻY�X�42��&}3�VDZ11�h

K,�8�CE������~5�`:n�o�$Cdj�-���3�	�!���Ա�/�C�z�z(`�d8��(Ig%���@jm�U�a<�;�0` 3�Ϡ5>QT˷n�a#h�S'� �Y�(�I���xKF�ЪX.u��*����̤@$��+(�K� ܵ�:��S�f0��!��t��p&�\���8���-��[hB�^�n���dC�(�\M3��l�FX�\3 ,5���*�2�;Nj,���p�ߑ���?��}�;�缀�f��,&�"��5 �M<l[�pΣ���Xب����E5����u��GΝ$YL��6��@���W�ʍ���s$5��NP�eޏ�ȅ��Q���Ytϟ �HN���o�>'��<�i:���d��?u4�`u���ko#) Ϝ��ʨw�n��´	��������#����CB�ӳ$BpH��uPW�0<h��t"��­�����,ǒ=��Q'�Ht��ۀ
J %,pY´t	����p�0#L��x��3�c��g\�|U�V�	lV��)�WD���L}<��0��#FƟj�R%�e&XmH%��U~�����s��kk�p7�ª�B���7䂄���A��T7;��HO �$K�<�*��d az�=d��چ;�E@�Re��܄�ǺbE�`%%�s�Cf�;�- d�
��a��<��G�3��;	B�4�-D���	��j�rE�V��wY�������ѯWZ ��6$`��h!�K���y�,�*�#�F�q�Cf}��4����b����V�E���x�X��nH,!�#�{u���{:�`���������4G�*���ī�w(��*��=�Я/� 2,�Q�͞<ee���}��sX�|��/S�3˵{�#{S����N=k������� "X��@���M��UNB�f���&��F8r�"�a���N�x�1P�aR�٬�qY:PX�X�(�]��vZ4%�Рz�����1��#�Ư-�C�]a���L�1xa�Q�W6`n"9	�� {�r�p�l$7����C�'�n0�TH��JG|�c2Oj���2š���FG_#�����\�K���^����|�҄�7@��}��=V�|>���fnm�2S� ]uY S���=�9E�+W��mr,��M��r_)^$V�
:�ˁZ���+Aݓ��G���w'l�5�N��NG�Q$���(N�[g��Nҍ�����+H�+լ���t�rzh�7�7]�+�Hٚp�p�*;��9�Ɖ������Y�qG}N��`�heq�������vŭH��@�(!�[���N��U����Tf~1n��#��
���v*�~���kb?�n�#aC�MPh�i��ō��k%o�Σ�/ꂄ�FW(C��@��}�I+C��~�#ubAn����}**!>T�[=I��r�+��EI1��i�c��C��5�"G����D0�`݀	�'NN�.Ͽ�FbOQ�8��$9qpb���:z^�	Y,1=TJ�s�o�����pb�� u��?�v�5�����ٞ�B�����$���X;A8�A#"|n�j/�ʯ�Q�+�u	��T��Z照E�(��^�\P\>j��F�%� �0Jى8[8���D�����m��Byh���,�4x��E������Vm��>�H�3&ռ_78\�
��]����� ��&N�i�ۖ"*��>D^a n[�<��4P����:g\�0l'��)��]�f�� �l�c7�&�X���<F�<>����DRʂ5���VhiՅ�CuZ�O:��~$&:)N�nr�:Wյ�j����M2/���'Q̙em�0O$�'z"Y !\��4 Ǭ��'\A��㑱-��`G5�RS�2����[��,׃�L�W���U*��ۓK2� �]�Y��f�Θ���u��@���kʱB��WE�&��p̐hn2!DW�K-�WZ�H�k�u ��f�����w��6��O57�F/�e��"R �+��΀�j�]�&n�H@ Thf6NP�O�X��w�w�sJ��KYe����T'�"zNA"�k,-�6v`eƉ�ȁI�pQYb@"$�Ql�<�������]XXǒ>�v�V�����	�=M��#:��j	�i��i/�r$��5��Z�{��'�к��.�u�, �����x�ca6!�0:b��Q�,�.9�Ƽ��*{��n�5r��CF4K+W!�e��:�(Vo~[���X��x�~X&�*� =�VI���p�����AQ!�uL~?Vy��ƞvX�<�no�¨D����w�ΗPN\�ه -��HE?H}�s@�]|�0���3�A��H	�qߛP���(3�qi	�b�M��M��>�;�I�:����R\*�]�����2��|��l�~e��-#֩��Tu4e���8�J�xN��mGִq1��|q@�V�>�_�-)��˞D��8���P��4��,T��Oy�i���B���N��B����/
M�z8+Hy���#я_�Δz�}m4�����F3�]�Ʋ��E�VQ8�άn�\s��s���JF{��芬529G�E�`?{�Sa��`F�D!�Ѫ�����/ i&�,�ZU�v�<��f����S=9e��K6���_���4���I���	D(�
�&�Cu�IP�X����E���OSz��@� �\�
��-�ʔ�9A8�guT�)R`�R:*�^b$7�%fD�άԼ�?�.�0�(C�hA�Ϳ`���4I����ZŨN#"Ii�e�S���\�hq���<��7K�0*��-W�|�؀�k�����j3rIڐj/cG:xO�,��`,O�\��6��YU#�¯'=x�u�G�����q(�jhSBI�hJ�2(�:�+�r�$�@���8y��r��c����^��!kR���J�	S,��d�m���]�X�mD�b���#JL<E�B2�6ȴ�+8���/�$�DMd�I�񒬼d8Dph i�~�:�1���	�H��{�Y7*V��uI?�"u�B"��4h{n�����"� ���M����Ȅ@Fki��,��L�\�N,.�2�R��K��u��S��:[i�O�a���h�x�qH�Y� k{"��C\��&�-�^؇<���_p2�-*z(�}��':aJk$Y�}ή�A9�/Ԋ=%� ��c{ W �IJ �I��-���x�8C	�h����b����0���)z!?3�LO�����Fç��ˉ$N_�M=%���TTCu�$��B8
g�N8IWi�p��X����jy�@V��'� �8�L�ʁ��Iq�i���%��q�"B�E�씹]�T#��זXf�<���;cq2�VRLp3U!�EYCj)�U���K���a�X��[�#�)�\��E3��I )8����{��^Pf�1c]=}�ݹ(8g$�U�=� �������{�̮�+<��6T9���;*wmf�����?"6,aa�dk~����e�&C
>�0��Z���o�M�y�%�H�d���V�0A-�̹#C5I8���? m���23w����[go�=u�pc���~N���y�C)���M�������6~@�&��*�_��Љ�����̿bn�hK�M   p�P��_1�s&�*tAK��;�%xJo\Ir�s��n}6<ҧ�j������H�ԲK�(��k�����R�
X*�!�^˭)��@���ɸV���A�<	Q��c��j�B��G�={4,3��<��o�TΒ���~]���ַ��������� �89^XG(���:vNbb!ºr��Z���Pn}����w��xUz	j`D�T� �XQ"��T:�Y}�_�=D���&��޻��񳼪r�4so����zweuY��'�b醙j,dn�b�l��F��|��zZ	ъ��X��94����ɘj&����C�elRZ��ct�b��}�G���[O,_�!���,����p8+�峱1F�PJ�fJ��1�������Oe ֞9�� �|`//�Ѵ�9�Z�ʶ�hGU>��m+l�h	^����9�,=�aU��3��)�6d'4{��`$�ݎ���8wX��;{o�Y^,�����?�R){�He���WB��) ˵B�{����~M�Djk����ԗ"g;jL�V�z�֑�i#���'�[������u� 0-Aɑ+Hb��� ����ѳD�WWߩ~�J��S��gNMʼ*�xh���V�$��eH�[�`����%_X<�Q���1��ǝ��e�S��
���� ã����)�)�f�/�ή<���J���UHz���LBj�$8����xT��v�өf�^W���4�%��G�f����T\�2Ѓ����۹��$�/`�w'YN1ezE��{��QJ{����𓛔��-2d��bG�!%��V��'��c���-R��.�IۧwC��J[���?�� K�8"���(�T<�}!�)ؓL�=�_������I/�� ����2pt����*1PJN	G���Z�q�ߩ�kv�m�o����v�J+5kj[�AQ*	�X�Ҁ1�b�?6E��L��)ƌ`6c��D)<@�+(F����^U����"�7mZ���M�� n=}I['�
�d���B�N��>1����z�%W˱������V��Mc}�����67r�D^j?>:����9@�v-��bf���mj��՛��g�k�����@�$���ڑ��h���^i���X�<�r*i�5��"��M�w���+���*+�Ý���)@ێ�?����ea$3]zC�}���h	������0������k��ջ��� �D}�@]
Ji�
�G�y�m��8VZZ�
v�",�r�"d�u�Bu3 ]N��B@���U��p��� s*����l�>��WQgU^}ĖB�:�v�)���.��yW0�n7�)��E�� � 5@ʿ��4v`�����2���Dp����� ��F�IƧPX[I�����x�dl�lA�,��U�(«i����A���̳,+5��9dW
�E�P�EP�U�WĈ;D)��l,��nS�EX}��aJ�ZJ��Tc�����\K`�3>HD�@��E����Ɂ�^)D����x!Zm���q�𞝈r8 �����B�nP�Z����,�I"��� I���U��<���N!KqB���SY�������� @��6<���E�� ��^�����VxM@�G�jq��9�āW}�{���,Yf�Vd{4X]ь;"
T�\�(*E���?-�@�s~�,V�����,9mGAn&��(�UEIY�����Y�vfԒ4
�|��oƅ����eIb8H��¢	�p�0����`�ZqKEoiƴ(#�[�P��ϗ��e��A���.� dʲz�����፞�3�%G����r�gǬ��bh�yt8�R���F�V<�
�@���En���Hĳ0�����Ywb�b��GMn5p�RC��dd4�Y��$B��rq.|n�K�/�2�
�� �8Y5��"�lV��d��{�s�B�0x>�� C�,a��K���1����
�����E��IEH_Nzg���.����b7�5f|�?m�^��n�d��b����W��q�v�(�Ω���1�V(�^;Y;bccQ%�@�u�fW�T;�v~O!��*^�lD1���!�TJ�~�� ��摗uN9 �+
^)�-��B8�S��T�0�����8��6SU�;y芟5!�a؝.x��@S�QV��L�-"
�

Ir	؜�,E�\N�șR�^r���Q,֤�JJ%,Ui`�8���
fX=�.� VMi�Ç���w�m1h�aܰ����1���84QB�Chz�c��Ŵ���K�GBl|~�%�� wUv��7�_v`���3U� �a@��E�
��,4���)UY��[�%������%���w۟�S�F4��d�1��w/~>�°&!ʯ�)�y/��T�W$��!�;��l�����=����x#*D;p��l�{
�WLA��V<��N<vo\9*�������n'���m�j\)�D3�-�J�r�0fLu�C�euWM	q�D�B��Îe���t�M⾐s ���()B��_Ʌ�����`��u�~@v�p�F�8?���	����F��Jl��u_������ϻ�骓X�t�
7�M�iYb�?������a�kϠq2��$D�!��� �}�dWn���t���7�Ѩ�y����E;�y��EeK�"F����|&�N��'�2��0C��fY��B �P�����X�����jX��wtz�.8�砟���Q�6%(C�H�F�M��1"�ŅP����80��4|5�-N�00��5�v4�W�Zj+|�� ��}���Z�g������ı"	~���@$(��{�(^{�-Z��ؑ�����K$���3d�cd����6#����i��倡/<��7CF|��X4m�Þ�A�xb�WP�D���O�6h|+��W(�p�՗�⦚@�^�#�H��CŊNp�
�'�%�x�ջ�y/��;+� �ŏ����V��	�!W�A�D'>x;����a�����-&VI�S[%v��b�b6� �,�.aE>Kgc�,c��A�_��o��8���K8��,�O���CX>�N����1	I�����������l�j���д��7ǰৃ��*�X �6IE���x�#��>s/�+�jg���شu?gb�,x�n��q���
bB-���D�1��Ag|�u:f~���6�˝+����ps�
��A��1�B-L|�l�y��	��#F.D�\�A0�������hy0x�R��p�Y�:��l$�|���{�ɗ�h�AԬV	s�ނ�Na��D�D���[�)(�e�II�X�p�ˋ�T�I1�s�B��m��,LO1�m��Wy$���ހ�cּťf���.��d�h3�q�DMg�J��N3���B�=���"��Cg� Uv�A��q/݅� P�$8�X0a�/ظ�(��ZX+�Ч���vR�ɦ)�/4��y*w��O��~���20k�T����6��H�y�� � o���G>ޜ�5�5o��g�`��?�L;ܼNA�uQ�tޙ�֦y`�;�Ψ��(;_~�	�v�+>��g�ʨ�Q5	��\���Y	7��wc�̧���6��\����~�;mʅu�GdN!r
��*�����e��ja�;�Κ9�*�"�f{
��L�OC�|����g��w�|sؽW̕�%�f�hz3�o�f�"��Ҋ��:Q�H�Xr)�E�X>�$��S�!��u��T0aP#��t?��v5���3a�a`�K�UD�_�hs��5���H
��,�ۇD!���y<=�g�~9�.�ۛ��E���' �Ն3g2�v2�>�Ʒ7��N���Ե��ޕ+�G�
���M7e5���Mj.?mZ4Ľw�@�x�D�ikp #��tB�$�g��V��^��
�r����[��Q/^���I���������Q
�x���P<���STMoVә݁��~����D3;M	>���:� D]a=G��L�&����o�r���`~<K���-�|7Hc�L,�W�k�`�#
���A�M��qmp����o`�������8�)>\r�mގ�BZ�����������-G��*2����>�t�����0���r.�!���kÞ��{�v�>��V�t��We@�B�T�F]�D�֩�W���7�bO����+p}���5�����2�(X�~�"�Џ�n����S�u��Wf���=��7��}�3�Z�U��)D�X�%����M�xuc}�? ��o��>�qp:y���)�JYZ".�j�X�~0�μb�ӹ0Av<�6Xc�S<9�V��בD=��P8}ʨ{��z���c�r%��2��f{F��Q ��Ϻ�ؘ�O���a����1��� ��q[��i��?=�����dx�{�oEy��>�Wۍ��  �D�5zMrb,�'1���!��bb,`T��(��Q��J�}o�m�5�f����f1�lr���{��/?vYk��{�Sښp��Ǡ[W��ѯ��աP�H$��=PC���\`!�t�2�b̩G��6�+_��uM�z퉨��z�ch�I4�X��-z�ի���sg��e�������b��f�Y�q����n}7�ѬőN7�[}5�LNf���d���٘�����3zcƓ�1��9��H�����8�'&�p�;��"�}���w���,��s���و�yD��lT�
 Huv
A�qw$m��{(dp��mb�)�V+J���9l���g&�܁����RVo�ō��"]KS`����pbpCj�h0ۖ��~�ukC\pǟ���Ǟ�\}����u���"�t���ڽ�\8�	�>�U$�	���������c�1�� �M�vܾ��Y�_>�M���>�L��� ᷼��2�2��ѳ��Z�i�/�-¡������'~�W��k�
خ:����%���X�`Z�w�Ǳ���}/���]�Љ�s����Of����������|�5�/�L;�j�����`�7i���f�8D�)�k7��+�}�1*bs�Vj>%ĢP��#S��'	XKo��afM���ч�{�ɟ�_�^�#h߷��A���CJqF1�Je��(�Zгk0ᢃ�ry�_�0m����G�\����S��bA��w$v����N39�j��f7`�I����ѵ�Ud}`}+�����ݹ˰^�AU2�[���p�	?�N;*��������}
�]�~;����{	���mo����c�	;�Gf�/��G�����L�:��ޛ�O��v��S͆�p�ч��ú�*4n ���	��fu7�;ءg~}t?<��\|�,#�	a9/�	�.�궫�}#\A�`���B�sS�E[�& �H���JIP�m���`l�v߸M�z��^��-%
$j-�R~{#�����:#W���,�N99�M^s��$�V~��c�S�(����Ba�n9�B!��]%����L��B��j�Վ�ֶFxe6+� ��Ч_����-L�d��e8��ݽ+��V��oB}C'�c	��[��Z�e�䠐P��A�J�V�mCn�h�&���_��J����:\e��",听�C{فG�	�w,Q PmG��E���A��p��X"H��E#z�J ҜiT���d���ɷ�:��ߝ��wf���mM��H��ٔ�*�3E��@�z/�4�vL�ep#�74��H�P�\�^��"րnZ(�J�c����h!�%O����8�b	�W���V�%�h��ajUx�e�ښb���2m>���t3&���Dܹҏ���X�d;��x9�c&JtR��(����F�YJK�P�G:��lG��!���x�$�fR�|�ݲ���	��	����Qj�p����'��L-E�dmR�$U�n��1���1&�ҁ���>���9�����y�d��$-�N�+'acȴt��dWA�-�mn����
3���G6�!�Ƅ��#l(�uUӰ'ס�x��v�|*|�Y�ܶQ�J�S�6�@��]O�4x��\�\l���<�I�7��䁍�z�dP`K��""�<Kn<�<bF�ؒ���U:���(�]L��T*�#�E�"�� �]S^�	�� �u<(� 33e�Q*�?C�1Q�d[M�s���!�������7�CH~��e"��7آ	-����W�oƶI�-��!��u��x>�)�f����6TgMԷ�	9I�o���p=f� It���/�1��K�G�[3\yR��!�nh0��O~��9��Z䒭X,J��m0����.�E�%�տ����!,g�f��R�@��-@gG�qHt���'�uHPY'��Qd�P���E�;���|^f�cJj%�M��tb��N�,��QN�^�ȖCՂF�1�kW���c|��h�j�(R���K%��ǶL�t״b(]xAI���'���Ϫ��L�$�.�\oe1Z�IV@Wz�P��u�✘|�i(���h+�$C9�	![y��W��1C�AQX~Y�wT[�ZaHU�DL�e'��t����d�"D@6>Qi$�9���Ǫ7�D2[�Q"��V"�A�U2��䁂��#V����y
�<	�0p��3�U0c�eP	 ��ј�R!/*ER\:@�'˂K{�h+�u������|f&�|ɖk�)�>�_C/������!���	S�±SR"��v)'�1W�c�O&�-����8�����)�D&f_6�B�3����(���#H�g\1�q;�4e4��T !z\�.ȶ��ݾ��:L�$�/R�N�W*"��(�����tH\���ֶP��4D�e��W��u(�T��ĉ%%��R �%��c��]Au�A"��b�E�ku�ĥ
ZK�����\}+�C$j�F�at ;Y�t��/���FC�����nG�ן�~���Q�Z�+��. ��z b��5;���Ү*>�~A�V]?�=IU1�s\d�H�e���e�2���B�g�@	����6����L��;�z�=�tx������.���%[ذu9rm+�Y�����(R=?��J�Z���1��}7�2Pg�%C�l����X��2�f�`��T��mҷ%D�+�E���kuEu׾(���ld��I	�-�L��.A�V؊��M5��{������P0�P�g����ڜ9Њ�Q��,�
ꊆ(�_`�`����m��&��D��bB����R���>\h�*l��P�{ �e�%@Ls��rff��/�EˬH���ƀ(N�DgY�`x����]8=�����Ku�G�9W�e���p��b+��J����1P΋X�D��=����s�bS��?O���@1�������2�����S��/ zFv7`w�@c����z����8��?�4�1�W���G	�s�E�O!Ձ���$Y��I���f�E!�p��Opc���Q(�b�LԘEH%9J��1c|zǿ!cXAU�&|6����cp��=�d��|�vL1�\W���$V�g1v�8�<���?�F���ܷ�P��<�|�ƣ�g�8%�(f9єU|S8�=ޞw��{s�ԋ�q�Y�b]P���!08����8:mh�x���q�Ǡ�*�|�m%S���W��e#!�SO?�O�n�.GCeyƓp핑r$�"��,v����G�+�����{�$z=pᖋ0l���'^�����Q�E�Q��fɑ\��������gb�������
��I���S%-�G#k�����%M�v�c����T�� 4���cף)B�JIԇ-�=����5�*%��h-�u�E�`�Iا�g���b��y��ȼ�I���/�N��A��P�네3�����������1��?�� jw)�(k��m��%�$^�KL��"{��)�,��z��~�~V�}z9M8﷿��0bP��,�T�B�d&�1��'��7-���+����Z��.٤�N/�ӗ�Ð�&��ݱ�9��C�84NwI �4�\WP�0�x�Y��4���9��i>0��5u�$^Z>k^y��]/L�
�U�]���CA���j|2n�n*���.��H����2��C�ƽU��i�!l&#s��K�<ߚ���s}y5޻uι�D�kI��ܒ~ԨL813m�/�!�<�*�=a,�>��Df��������ܗ����0��?������JA554���o�|�<��d:������mH����t
۰���7��O��� �BG��XX��bP���G���K��㗗b}P'��m��˷�������0(���c����������%'�(=�׏���=�qH$�N��P4ѫ�����������a�%�����A��(��TU>�|>n��A�7�����#ű)]�(橮$��-iW?�cx��ؕlm`P���	W��O�A�v�
[�8�}��b��n��n�N=�bl�a���@ul��ٝ��r3
_��E3�Ľ���sr�^!�G�w��C�������ć^��LC#:��'�&�Ð�7�?V̺=�\z�)(�R�G�l��lT��-<��ۘ��~z�zW�%�a(PL��b�[�`P|.<�h��,J�{��x(�B�(�D�������c���E:H�d�����!j�,r�����'�����Y٥2�i$( k)�Y5�v��.ĵ�c�K�Z�f��y��F�
�CK2�nz��Ç.���}+F��U�o0{�8�̟���n�R��J0d�� _,�w#��N'�n�]���/���o=����.����U`�&&
ӌ�+���G�c�3��Yw�I�8�F2։K`�Κ�[�Əu�O9^�����nR�������k�t�p	��C��rXF������=�]��8�!Α��L�GG��G���'I\z����W%��Yh�(0�Y�	nM�An��X��$<0c<�0#T���^�v��̆i��}�?����h:�esVS��9ͷ�C7<t���;:[#���训�[�/A�6zVs���8��#��T�$�d\�m��9+����a��[�&8̒�@�'�d��g�c�돠W�ZQ���O����a���L�T��M�7�1�tkD��*�0c4|���h��%���E�n�-�uM����$%��A����v'��Xl(שVT�(߅��]w1���W����@)��g9P�!+.�Xt]l4�6]    IDATZ�G���=�d������	�*0���#��N��$!8w�]" 0��eőI�֬�2����"�r�g¢=�f��Q��#2�n�|�@���N�2��倷��ӈ8GC9"���'���7ջ��(������>���� �44��$c0�G�Mōl��z�����J�1����)��7�OF�{��K�
�*oL�����
)��j���������(��B�́[���/_�抗p����e�2��t�n�$�NSs
�W�ÂFk��߯G"�Q���-�d`�m������Nئ��BlM 5�RZ=p�$�����Y�A܇l� �=�Jl. %��g?W*r���#2Sƍ�2�ok�:�RcL��Y
������P�{u�D�^�\@��2u���y��w�ᱏW*;�$qL�����}/B�d5�$���u]��P�6,}{Z?z��6(�]`(�;Ճ7�1���h��Q�Ff���Z�c�;c'�K��!�٪(d���1[pc�����o���6�S.C[�V�y`�-�-x������
Ze�*�@^�� =��ɮ��kZp�3��ЩhM��zEށ�HW<X�>[S�B2��!c�K�A�o��Eӊ�� �E�/���t=n4�|�|5�C]�@mЪ2�_���xE�>c�I`�.�V/����tc`p���uT��X��T9JPhS�+Jn3d�o��p�a�?���Z�h�Dƽ���Z�a��b��|�8��\��v��.r#�IUk�������C�þ�C�슂�XJ,�J�+X��x��?�����f�!��F�k�1|�]x��T��pK�:�)_)V7k�.�:̾��ck����G�Qbjō�sN$%}tbYj/O�	�l��$1� �Wc���W��lW[T����Ӓ1����(ql��0m�?̞�k�#hһ�d�Na�Д��1mt�rX��$���� �m�K=u7A�T`��AWs�C���c$0Ȱ־؆%c�k:�H��'$AL.-�?�dZ��+K�/{<����U���E8p�uh��Q�و⁰]�`nn�_��������7�U3g
�W�0�V.o���ߏ�gޏb��pEԅŪjUU��L����%Ό��_�Y�������F��hYf��c_�b�fg���eH�t |���\�X��3��KX����%RXE��'��(�U���$�%�e��֎%o݃���_6Z�o)c��<J��NR'>Da�:������-6�O={)ӤӵHʜg�{�rM��xa�R<��2|�x�h�ȋ|�rT��@������Ϸ������\ps?�M�!V�FkW�1�ҩt�d�v 9z"��Y�$,����l�J:[C8����������|�΃�=�.<� 	���M�h���!�!����K��c+qȹ�Ь�6v[��6�翈�/܊�R���U���I��r ���&��L��
C�ƣZ�ہQ)>�gq��}��{�}\\��#z*0��c�o�c�D'���*��V�]���7���'W�a�eW�)c2ǨC�
��o�\�����G�dZk$$0�����}�Ԯp�}*cc`�(��O�1�&|8�5����'��Y`l�^!v��o��Q�Q}��c�;ӱK�s?y�L.��SGh%0���3�%0z���=�Dʄ�oC2F�(QNӢ�-���}����r~�!d�v���^�"5A��*��%�����*cl)0��І%o�������of=�]b���S��S��.���&Vn���-#�g�X���^�μ�F�ZLىs���$;�%,z�VL����ƈ�π�-�-����vu#.���{xc`���f<�X\	.�v�0|[`�;���E�?��x��r�hp���ܩ������Ģj�x�k<�\#�=��#�(Q`]���7����W�A�ƨ����/��ƚ��(r�ChO@��*���/+̐�f�(08����qS���?[|n���]"-�h�!����(����ͬ�%1眰?b�n�$ ���R���T��*O����ԂCϾ{��0�!���ƌq����I`DXN����5\|�r�	�"��� �U����c����jծ�WG��q�TsW���x�Q�nǏA͎Rn]�Ս6!d%����G��g����sc�*����yMܮFʽ�I4�����7�`���C���f��l\.�L8 �0w>�~9�A'AZ�vՐ�j�YƂ����g�boh��"x��U5�㢫H�.k�x���x��=�FlM��Kl�.]I-T`,~~n��<���;�!s	�j�F����hn*���f [����*��H��H�[�0�%wt0clu`���u˥���׮��
�D�@i���Φ
�@����	c�;��D��Q&G�z�Da���������̀p8�D���� �L����P���^8`��X��;aœ�������q�0�E����J5��X*:)�X(�}�tv��H�]a�`�� +�8u�,���ͺ(m��nQ�{8	"A��ϙ[9Qt=��8=!:�$o3؜@C����YX����(T f��m:x=��*��C�`uƐKF��[��U����&�Lc����P���1<�!���|�yԖV��)�����Ñ��Ќ�4�0D�����}�DJ1�`�̳Ǣ��Q��"<V�q��d>���.���OM��i7�*ge�,�]�����cq���LL������bu��0�sՈ�4b�<"�6`��5}�+Ǝ���%]�D%���2�MA4���<�����Ϯ�t�d�Ő/;���JҘ���(��Pn�n[���^@X���iZ�(�C�z'`�ð���G:��lR�}�cA�xi���c���&�8�%J|��.Ǽ�1X�eW$,�FW�>�N�]	Q�X_P,(����C����FW����/��'���iׇ�,S����1�D!���:�3�^��'\���{��ɹ,&wT�R�x+��WON���7���&Q�m|�Es������[31m�+8l��X�s���+�	��t�f��wr�?��7ހ�����7��6��$P٘��s�˜����[�5�����<�q�bէ/!\�
���2.��8
W[e��{ �F��W?���b�翇"���)nw	��׌`�{�������"�N����^�!���������и�<���06X=�JMXW�*2��i���d�E��[�]%����s-~w���>��0�O�N�-Sp��G^	?DU���`�IW��;�:���g���!��ފ���wb��7
�U��h2P	7��ƛo���z��=��t����Y6���d:�����B��R����:�nM�|Y��1L�Y��4��^��F�b�������ki4��+�_<�i׏j �°�
�Vf@9ЌLC�$�>�&^��{��9(�c�-M��@��_��z�VL��F$��rW"Z>r"I�$�S@��͝����C.{��9��_!��5�%�a�n(.���YcL��#r�[�J�x��
sf܌���$O'1���Җ��%��ō 邇sG^��']��n0�<i�-�Z�Q����]�}�nL�~���hW�5*�c���)+���x=��>���]ap�	��j��Q�7���h]��p�h$l�|^p����@��`Oa"``<�>X����^�f�q�\� �]#��x���9o�<�\{�Ŝ�tX1d�98���� �g������
{��TC�E�s%�"��E�1wL�Ն+�!&��`��D}J+-`���q��ǰ��I�$���hZ�0�Wծ�����gv�͗oY�sk�:�NF>��z��ȁ8���D�F7
��ȵ-�����$�<�Jl�eH���+��LS.\��
2(�x�w30�c��K��z��2�$*q�iZxc�'x�Y8�;�����?d��P����P���/x7����F�����`ծ�M�l���䳘��Z�s��h	����h��^��z��(~����r�6�P"�1���J98Ҷ�¾��ԛxc���q6�<e+!�L�N��O�[��>:�M�*��R�n�w����Z���/>����u�DdR��Xr�P�&�3c`H�U��]I4��Q�52��׺M��;��z�B�{��r�>��
�F�1�k��/F����(��7����OF;r+>��Oލߏ�f9#P>���� 
1z=��{}�'��9�;���e��� �8t��zvγhZ�.��L� �`(-�1p�LN�3�^���Vf1��ñ���G$��47���_�	w�L\s���͍�M��x2&�~>��GJ#q'	����xk~��rZ�*xvJ�	nbƬ
3pW���L���nAJ��&��h\��|���O>��w=�C/���ZvJ
Ve[�D�,,�EeC��H|�ٻƏ�ѹg������?P�ٚ� ��m�g�4/�P��\�7��*��h�����w�����"����5��kHy�W~��OL�,@9A�0�s�����
�ͦt�{�~9�5ZY���PS�;�e�9����y�)�
�z\�i*쳍>W��ό������3�E�������O��Âw_D~�Ӏ������Y#�+�wJ>k�w���Yhu�(�D��`��D�5_�GJ,>�AQ�d�.�]�l�M�����7!��A�>?$mG���䐋-�V���W�(��_�PfI1�*1']5"�Q �ݪ�!w�SP�����p�6X�Cw�$C+�JǮD�v��m��I&�Id�:x�S#=O�O��LCa���3(�����Př:��� $7��L:-w�'��������H��ڡ��dh&��� �K�X�{ ���q� cA�A��,�X��6Ӣ��+߈r�(礫���RS���&
�r��%��V�u������T8��3�>F�Av%�]ݚ�PMlK��s\�E�vQq��"G4?�c��Z93%�����dh�	�D:�t!��%�>DBHɂ��Z
�h,�(g����F�r�f4Zbmn�'{J\��4	�ȅ��
�h9+%�9&��X�j�S�G�\D�C�D�R�VY��5���j�*�[�(MPC�5��,^U1�4�*���G�Q��5=JF��O��K���HoDv����F����N�����KYT)Zn��ۡ��QZ���O��dq�)T�@���``�W�GR�\`ZaF�!'KD2�7�!��vI�óU<\I�*?4:-Ẁ%EYC��5��*Spefǉ!� �d
�� s��nW���Vv&JF��7C��L��>8�si���wM�2�4آ����
��+�X4VG&�Id�DEHyK��B_�B�b�A�N�&|<���qc�lή�a�8N��LJ�GE֖�O8J∁$fp*�q��񆋰�����	�;(F�h����E�1A?�5��Qe&U�(?CYw30x+6mJ���r+��H9Ϡ���d��qE��d@�x�"'�x�����H�Ӕh
	?�A�h�G?V>,q���SX�>W0��uTΚ�<�"j���=l�"J1�;"Pi��cgS`��K��e�q�O�9�w����羇r��^�p���E���+�n��7F��se,���QN�܍��<�B�r� ଟ�H\�g��cD�YX���� �y3U`��T�/t��&�b�RA+�e�j����<���Zo���yLX�|<.D[e�d�<�|���`�̈M�q�������J�F�|VTT�#Z���f��k,�~����U�%�kb���_��F�0�Y�D�v'�:Jd���?0$��jW���RW��M�'ʶ|���QGwm'���L))FUᤊS>J�J�C9�#�J��O�T]��U}Q+N��h��Ŧ��V���C*GG�1(���a�5��H��V��,<�� r��p�$yE�"_�~��<�f/Z�c_�1R	�cS��UQ-���QD}~n����/T楊�P��7�j5_��m�*>͍��%0�]��0o�|*K�
kL.Nt!7��Q�D\L�F��H-��,�<~ʏ����0��i���>E�x��,R�Qe����Ճ�o��0��]P*�D��v�v�8:�虁�T&=<�:\I&(}�YI%}Nf
�xx|H���[&��F+1:�YC*�Q�I�-�3k ��{��M���T���Mq7EƔ��*G�a�{D�I�ԋ�Ht�5�>�L��2~�k�i�fy���_���$z� Fda%$ y��gy�� WD@9R"־ �&�|�����B.x�RE���UlO�K��At�J9e>i��������.���{�*y�6�n\Ή�w���@��ZW܊����}��V�P}$�I^f&Փ�5��B6�Fbv$�������fS�j,�U sr��ḷ@�����"e�����ˢS�g�L�U�*���Z�!hפ���x�'���o"�m�#	��ƿ���N�W7����sjE�&�6�+ ��_Ԏ�8�����eJ��w!�	Ӷ�泈9Ԩ����F����rY%���!G��g.<7�H>�eU��p�u���:M��d�Q����S�CPwӎǐ)����e����ԓĖ��\����J�@��N"��Fw�جZc��0�(����%�^�Ϩے���Q�]�Q�ߩ ��3T'�^�����p��ZLJ�D�+����~��ˎ� Gn���:z	E������)�;��<0�4"����e�w��=�PB])�����/�p�У�gY	����ؘ+�q��P#E'���E*���2��)����Z?�[1�G�"�T��ȕJ(���;�QA���$� vٓ��O���,��*�b�Y������ి�WZ�ddN���rQ���ř��9Q��/X�Yp��y��ٕZf������k�����W
08�|)�):P<�|T�.�&l~��e,����}�y�:t�ɟw c�$�I���r��(zE��h��PcI��>)�Y ��E8�����l�[�s#6��b>+j8��EN�"pRhn/"��H�yT[�ީ�Y�n�RI�VR���� ��D�4��"h]���!i���e_d�S19��t�o%�C=z��rU�0Ljp� �����D|U�ln� �K�А��r������m�U��j������P����t+F�(q�e��P��ކOo?==����)�30�L�q�ЋT`�G��,ʬ���վeb������m�ߦ~����5��D��jt�H��֮Z�uO�n������) Ā ��/��^�\��;��mR3p�W���� ����ߧ�~���g����? ^���m	��~:����g'���=��hhk�@=�a���3b�Ӊ��bI����{�V�dQ(f�b�����؄��
�$ߑ?W6V;���S>����IU��to|�2 �!t�<ЬYX�q�������a�n�h�s�8��-�ŷ���wJ`���<�̟�}��?�;�E\s�0�n�I4���E�[����?c82f-��.C�����᧣*��!�=����m����Ћ�AZ�F,,�����нk�,�x\P��ؒ�0��I���@�'bz�O']�a瞈���F�Ǜ@�=��6�K�n�Cp�1Hl��}GIOS����X�(ss�|ci�r�Hؾ���~�Ѯ���Yx�F^ ��TZ�ʤwk����r:.��P󞲡8V&*�]TQ�4\ɦ�N}ae�0kҘ�)��w��n!0=r���7F,Z�t���q|�.~M�&c�u� ȳk�P`�Ӱ��9��F_�Ç_�l�;��E�;�q��Q*)�5�I���_���u9\5�&0�jd���i|t�Y���PW�I::'��J���>���$h�,���]�\w�Ht��M�b�]�_b��%�c�� �Ͼ�Z5���^JY�F��m����o<�`��$������b.�,�D��ǯ�АB3*Z��T��D���Qc\v-���<�Ja��F��^����)�H _n    IDAT��r`L��5���>A2�Fw*��qѡ4�,¦�X��͘���ÆǳMv:V�p��q8�?�9�-K���`�b2�v�w�"eؖ�ōy���Sq��k��o@����[~��:]z�Tn��}�]Ӏߎ��G��t��Pk���� C@��q���SC� di�(]�����.����D�Aڬ���E~ ��5���%T�!�~�6r+���N{��������R�t)�#E���������V�r!Tn��a5_2�ć@=M�\u�����-���F����愑�S�{�g�����.�7md��Hī��K��c���q����2� N��� vqc��D2�hKl��_�p��I��9���N,��0e�p�Tr�MXo�@�܌�������.]�t3��Db�,�4g��=~<���V����N�M�G�.�jmz�5�� ��8{�x:�7(��mV'��!�r¶��J
��KRp�9|3�֭��CQ"�?g7#�P����;	�������h��uߴ�Wˍ��7����۰��u(��%> l�"��D��a��/��g��]�O?f���>i�w%��y���G]��!�!��'5�$P�*���UBn�L�|�6<x��02=A���t��l��އ�-�Ѽ�+�߹��*O)�8+U�|����a�~�$6��	��[���ᦫ���[7�+(�H��bX1\x���w��ж��b��y6n�r(���	ߧ1�����A1���+nĮ�ׯ���j�2�L8�kg"�5U(b�ϡв;>.�n���Y�W��+���X<���+�Ҏ�,�Xl��L��r���"�Y�f��?F�b�YW2l����n���-v%*0���!N�zԉ���q]"A��0���oc��ɸ��+��-]�h�h)��e�q��p���b�����c�_oÌG���#�K%MGm"�EkҸ��;p�W�X�z~>��t�t݅���C2'��o���bI�2l�����:��bָ���G��s��� ��I�z�F\�}~zܮ��uF.�e6!$��إ5�c��O!�Ҍ��OKD��h�(��j�*���\���d
���o���h��� Q�r����2w&�\�O+�O�Ƞ}��h��)�I��w�<�}��1z���.>�}��]��z�A$��q�H�W��Ϟ�.*2J���N�c<�i�c�U7��F���B�j)>Ǐ��,Kj�`�r	�(����f�q�yi�q����O#ѩKW��p���i� �sɕr��ﳏ�-�<�R�r�p��7.#���������O|�Q0z�\�rNg���'��U�6�a��#�܂���	\����Z�݋�W�[�"��ʪ��q+�cK��nį�*"�c�U�SE��V8�72Ȭ���9�c��k7|�?���I���rƘ��މFԋ�,�Ǧ�"�r�x��JM�.��#��[P�P,p���C[��ܯ��?%��r�V|��A�vqF��[HB|��$v�y$7�(|��k�uie���+kh��;}���;�K������y��CUu��Q�.�:C<��y�=���Z]_R�������wV��'̰��ȥS]����E�����%�F��j,�\"��R�������޶�����T�&E�BU�wZ��d`�H��ȭ~k�|�A�ƉM��m��Ʊ�w�	�;�1�~75r:�|������ yq�!��2c�+^X��S� ��a`O��� ����^�h@f���*rT�*�����������Wym��y�op����g��9�Y��O��M:��[�Z���E�^��lK�r
z�,��U�R䏋�����Q��i��ŕt���
�韼8W�Qo@$u����|���H�iV����nD���ĳ�&�u���{�{��3G���>L�F���y|���(~�*Pj�11��!��Ӱi_�`#��T���-�~$��L8�ݨ�Z�ԱPR���M�'��'�X��^v���d_��~������y2�R�sz��w<���*4y5HF�'ї�3c00x����g(j��J`Tgj$��Ѱٗo�P��e��E����^S�6z�S0����QQ��MT�mȯ~Ec�97#n���1��1e�#�9���O��A��ڰ+ߞ�?[U,Tn�T=j��p��1Me�
Eo�����4��=A��Wc��z�	eSs$�V,�D�5V󏲌���B�ΫG�lu�������5?G�
:g��n:��Gl
��<���D_G}؎��@������V�By?ɵvEZR�6��Q[l�eC�yM�Q;r�ȕ�����A2�����&�FJ�^Ɗ/?��a��1C̾�ܶ;o}����E�����!QX���ߏ5��EP���iM��$�@��ʲ�B*7K	H�/b�*�XL���h���h-�D�1sk+.F�d�O�	������E�1�����U�4A����@��� �_�ɒ��A�09J*�d����5��ϐ�E5�ڕT��Y9"3G*Ҳ��M7D��:rR�����_�
C��b�QGö��$r<ʨF��D�I7=���hcq��j��ȶ���ӑ�[P\�*V~�)vv�pwgO�6��Qm�]�z�?;����s�9J�%袷c��w������J�<*�Y�������Xe���:z��#�n��Q2Q��+�o}��n�6
�Ejn������=O�f��@����y�}������������<
%t��a�p���"7�j|^q�L	��M�TA��(�@(��O�Q,{����d09�Y�T�������!(;ΐ+�2}1���.j�k�Q*����]Wl?.�X+;J�Q�GU��.i�"��-���s�~�8�u�(�)�F��vu�O�쬋�v�᷋!
U��X��d4}� _Ā~c���&����6\Q`D ���S�CJUc�������lt�AfxCd���lW��d�=���D w�C��r�(�[ø@�C%�O{��Eo܄���hZ�ɺ8R5�ZĬ�̅ׯ@�ϡK���)heq-@�m��M�Wա�~�~��W."nSۣ���Ĝ�VJ���!�������wb�"a�!��]	��î��������#�=�-0: ZDj&���.��$� LG��Am*���q�b�N]�u�V!$.��G6ׂ�_D�>}Pv������epةK7؉*�3��H!�H+�ǆ�b'KvB5�g��e̱���H`�}�Ň�s�o���Q��|[`t<c���bNc�%e�+-&Qd6t��$@�Z��������%�;%�HQ�\C�i���	͙ft���U-{�L����X5R��a�q�n ǈڬض��ص=`�ꐰ���,il��2ƶ����EdbQ�J,#0���D��Cw������"��:��>GU�ӱ�f�R�.Q�9��T�����k_J<��g�y�X��ֵrĕ2^�K<U��E�L9'lE`�O�e�!g�~ʗ�2��Vc��͔9��3�	����ۑ͵�h�[�ż7���K�h\���z����~{b�;!,瑬������,�[odJ@]�t0�^��b��ڶe�'�5�K�2�$ I[� � ]�t���X`L���qC/���m5FGj��<�E�̒#@!�Ќ\a�����n@��yX7�E��i��ð��H8:���!t��HR RH��X�f-&M��Oޞ�Ԡ�ѵ��j5XղN�
U��H�k�20ȋX����-0Tq�q��NWB7���(#�s��mhA3��%�
��ڴޒ/D���}1��Y��t�2��k�����r��q7�/~Hv�vA��.Ы�Qݝ;���Ȓs
>�f%�q����e�m�gǋO.����Lő˷�n��Bz����n��/�Ev���i���'�
z�ҥO?���Ԇ6<�G2a�-�ʮ��;'ބ��yI��v�%�k֖�������+Jb�ǀ�ʐ�FB��hJH��]|n��{��� ���|#�$��!��)�cݢYh�`�;dw|��,����pvۡ�?�ڮp�	����T�
�n��?�$vؾR�:|>ov�7�7����a��G�h�@10�1������Q񹱘�B`�5~���uҜm���T|���	
�X�~B��TM
u5lw=�~�~@[#׎�{�C*Y��m/u,Y�5vݥ?�|��;�X,�;n��=�,RH�-��yTW�b��ň�vG[����T�G��i}�X-��pI�)nޕ(��p�o��]��G�F��j�ge^�Ѻ�t�3�塃1�曰]����j`��siT�m̝?��&M��rp�mwcƣO���3�V�/+ee��_�#~zjz����?�����������I`P��(|%I��%0��ķ��ಋ�������V��^�����57��Q��in��ӧ��v���HC�|�,�f.~pȁ�a���6�A���V<7���\Ĭ �����W�m(���OD��' ^������D���@qy�T���1��Vo��X�+=�G"��^3kg?���<�r	5	wO������N�z������KX��B���ؿ� �KG�/�tt,\����wO��{�~�����p��GB�h"@Ae��E������Ə>d�5ƶ��x`��:a��Cqo=V}�:���b��W��n��X2Ҿs��x��ѣWOh�rՏ��4��B/�Ìk�X�p!v8wO�S���୆�_zS&>��G�����^#��[�%���m��q����U2��p�lW��liٴ]�pj�N�
��2Bz�S���Q��aeW`��᷿����XP��a� ��q�ģ�>���	a����!�l���F�f�B��q�u�4�$R(�6(�����e0�������Ъu������U'W�1�*�@b;h ��G����[F�ő�^�Px���j-��x��G"��.>�z^��L[+�f�&���r��FM����^���g��]+�懯�	R��*�m���ǟG���#��R��8�X�r%z����M'\����Q*�D�xyc�=�|�8�8��;�A,=�T���j�AJ�	P�N����0=jpu,0�L{�ء����H��fx��<�Za/DÇW.��ϡ�����FQhCJˢ�q��S��:)GC>O��j�	�x��'0a���ڥ'�H ���͵��@{.��+W��_��]�r��N�8�l3庐�}�I{8���Q��1�[���U�db�*h�B�3�-*G�1�߄��,����,0HhA�=~��Q����S��tX����CY��y�V$�~�N8nW;�(���P%aHc���3q��Qߩ�D|�t�@L)_D"V/��_-���O�F�w�L;H.��6Z�"�l����n�8�0�Bہ%��}�H��|Z��f0����m��OP���y-?��~��D�n��$v�bl���X>���]�{o���&��ke��ʛ���?^�xʑ����#�+#��(��T��r��`���8�����s��%?@��{�K�>�8����5B�jS���QW���1���a�؏'�߱��=�=v̙#�=��(Q��{�Rr�)W�����ĳ*$�:(�tۑ^�!�~����}��-$�$f�������Zt�^��rG�������跣�a�FOk�҅M8o�i8��(��$F\5�8�~����6<�23���ZEE``���u�l�`>�;c�8�h�P�\�IA`�!R�
}]
t8�!SJ����k��_��d�r9�{W|��,\~����E}������NҶc�U��k���w�{��B���I�
� �+�b����8���p��g`]&��:����{�r,�2�vĲd,`�HuY�%��m��]��� ��A�;Օ�S`N�V\��22�Pη�q]��6-��~�4���#q���ѥ�u��#T%Y5�<�����ѩ7.9
󾚋;@�/H+L%�l:�5+��1c��1�'~]�9�H%��RH:5���h�
泂���w	�=*>�e��g�
J��t%�(a`�e��u6�'i�C�
i���
��кA)��d'����2������Q@���I��!��a��F�iL{�>���&��=࢑���/�`��v�C�PSǒ���u�n?<Zjg�M�����������V�0�-��7^|���S�}��]��N��9}�Y�2���n��V�;�'X�Q*`��X��X�L$�<J�s���;�`=�î���Ʀh-��࣏��Gg�b1�Z2�IT�m��W'au�Zlק�N6��Wd��G�.G��.��d�D	1xAA)�TT���d&"
;¹�-0��v�bJFd��� ќ��G`�f�+ۈ;&� �}V�{������4����+��@�����|Q�3J���I����,D�.�L{�k�d/��o�E�a��M��(+oڍ\0����C�S.����Y�F��\!)�%EAS�#�+m�����(���ˮ�QhDz�B俞+,> �g܃~�C!�G�U�l[;�S4��3����1삑X�p`uj��ǀ��%�h�+��U���f�N�� �[�wQ�����dE8j�P���Z�m!0�T,v�k_�Ppې).B�!Z�Y[�̪�X�����y眂�T́S�P.`;:��툧��vsXٴ�~_�nB�� x8�2y��6���n��B���6�]��١��������1Ó��2n��u*�l�9�SB*GG�U|n�+��E�L�$	�U�as�ihI�E[q9KC�n;A+���䱦1�� \C^�0{����llhX�҂�\y�qe���>���]Q�Q�Kؐ��"i��.]�"�̒XT(�f����&��VsW+�Q�v<0�+��+��E[��h:ׂl�
;�e��)Z�#,� �~|/-���6�X�0ӪtA�����F�^�D����Э��ր����iȕ��PLCגH�I��d��|^��
G��#c���Z����
�o���f�^�����@;j{ht.2�۾ȱ�c¥�L�J��mH��D��Z��8VI<泅"z��߷�[6
���7ÉU!����T���D6���DcLi&�"_-v'�B`�9�#RKӨ|�K���۽=b�+�v�7�9���T���*�"U���
�S��x"���FÅM�����~j��6�AP2���O�B�?yM�v?�Z�Aw �MP���3��110Zڰ�?�*�Q)�"��)4/5�Q)�b#�klx����;���v�hȣ{��0�N(�<z���s}t��Kp§VƲ��E��o��Q(�g�$Cp�B������9�)�U_���}�U��\}��8tQ)bP{ID��D����E# �t�b/4iV�I�����X��Ac56l�H?e�U_�����A�9ƛ���Խ�����o�D*4�����pp��;>[�s���ɬd��=�|��aL������Z'�F
��gغ�Q|��@�$p��t@�Z������lJ{�$�o�`P�l��P�l��'�B/:&��2-2��kCiᣳD[AFGb��o9`E��=����M]T��),��;u���g_���>�=EjbP���o��j-�w��0�[r�9�L�Q],#J��-����!����4GQ ���b	��B�RSW+�B8g�l�Z��ܹ3L3%FB�%~��i�02)�LR(%�wa۴ќ/���R2��:\TY6�n1��(}��%���kW�8�8���o�Ըtᴣ�H2���>y��e؈��2�I���O���~�[Q�4O��	q�h�)�+ތ�C�,������$�P�QsT�D$�P\\�pMPuȐV���S�9�����C5/�s�-�'R9��I��0ۨ553v3bR뛰z�cF,�{��vJ�7�XDb%������5���u"�I3T�E-ơ�_q�B٘���Js�ZE����AnڼA���:����P��#�!)�lK�hD
���ɩ�}!Zr    IDATj"��ޅak(� ���ס�<�v����F�c/!����7p��kP�ұr�؆�g�G�ye�<|�2��4B=�<������'� ��,4r���ي�Fi�JH��b��%>Q�{�LD��\C{��Nhs��n��NQ��X�r�[��1�\V�%���ka�E�b�'�iH�%��d9�>Ǎ^�sRB.���dV�#4��x�韢����	��nC�bT����Cc;�,�:c2�XS+!0QR��c���Ii�567H~��f�/"b���J�4j�E}�!2T����F�q��Q	A�sX�z��'��ٹ�lh��Z��nM?�yZ�?�������n���x����\0���#.|��y�`�d~��76i�1<T?ŧ�����X��3�C�V\,�Z�J�J֜�[�3W`Ř{� H�UIO*��Q�$HH��,A�����4ũe���:�*�'�YʑV���,v�s���p�5ȥ�F�q�/�7��I�T�7�ݧI�ք�π���0���Ȕ�"� �7�2!������	�u�X�3YqJl��V����6��L���s���Qc��7�q�K�2�48�V�4n��:���S�d�l}g4�}	��~�.�]:����?jX>��^z����{9�ҩ~;x�
1.�v�6c��?��g)Z�L�l;����u"���w����X��I�.Z,L�b�Bj�^��d&I�`�F�4a����Z����\1���Dah�G����D�����%�6�>�c��3М��J��[�y��4s�&��_�Za�%D��8��r�bK��bPI�Ee�C]���X�'?�&�y?�kN8@���0	��g��(|�7����'����"�����~=�{`%:����7�v�[8�2
5c�	�o��g�P<��M�بu����h�[x���h��v���J?���PY�#q	��Ɯ�%E�J�j�>:�.�.c/@"!�R��"��1�o�y�B�R��\/'�=���>�y���͘N�3����<�*lF���N���n�ZcU�2�A߃�*��GEf�al�S��]�*�`1A�B�)wV��$���/f࣠�R<j�J�ÒԆ�S��N���b��	�ϛ��	Җ
U|[�m��`������q��}kW����@mFów�m�a,}������Ѝ2RQ��#���PD�[? 6��C���,d�<����%��5��kV�԰��.�?��E�+�NW�X,�6-4=|��&T�7�ȁN��G�c�^]PW�UR��:	]�g�a�+o �Wo�U]�IYBF������Z%�#�Ym����kk��� ��л�~'��f���	�p8 υ�j���EMW��|T�5_��";�:�ݫ�nb���@�$��*���B���$��T�(8� �9���C�ք�����3�ǡ�:I��n��,�nC���}�p��*�}�uq�lT�����x֞=Ʋ?�FOX���/_&��je�Z	�pa��3"�׿�w���͞�Դ$l%��i��E�dS#���f���S���5����a�U��0(�+�S�j�ç[��>uN�t5�tG�yr�T,Zp�w��iQZ�q]rz�6�N���}6����񻅓1�4�ثtS����*\�pp�sp�)g��r��.؊p���a�O��6��w��
[����S�#�D�DAY����P-V|�(?��
 ��nI>U(�5p�����bOĤ&,�P�0$f4�]e�%+_�߆N�Vl�`%��9�׌������6WF*��>��^_�A��$�}�s\������|��vH>������4��G_~���
^	Y;�XD3D�����_nŃ�_�BQ1�f,�b���m.��q3N�trF-�������Λ-(���g����?ؐ���ޅ�_~���T���E�1o�$t�I#�Pq�D�lW����&_�#�}>r]C�����K0�dt�Tˡ��&�ob��M���N85}��Mn�Q%��|"�闔G0,9���(�K|���1ĵK�h�Q0e���p���H�n�H�͗C�*dZBHk�XT�_W�=t�Aa�:h��H�p��Ǣs]=r�2�ٯP�:�G��g�J|��5�q2v��n۰t�{6��~��.7�_w�FI�D�M3��<�a�5���g���y�����Y[��r�J�̽�;�Z4uȯ���~�hDl�H#)%Ib���ֺm��{pԴ�تף�^ċ7]��7�E����x�#]�@Oa��Y�u�w��_J�X}�E�oҵ[g��s���=�U�Kf-�~������{Ҍ��+��bpfE&q�
���5O��-[��E�D'����+Sb�J�a�e��l]���b|�{�y�'2Vb���f��H ��BQ�yL����	6��'�|ad`�����ա���oF������8h�I�_����ƍ�8��Eبգ�
�vP�-�P�|��>�w�0�Q+ՉC�t���j����믽�\v��m��-�_�1n�5J�V6l�#�"����<���n3mևu�E3^�w���.���$&�R�t���ԫ�����A���Î�xc�EXx�t��M�C]��G"�9��%8�ĳ��<
[�l�c��Z�J}��N�#<�[֭E�#� ��3��Vj��<��	�+��V��Vd�w�w�{�%C���B�t��;�e=�7�c6M�m�nwjPpT�>y���M^$t�/�~y��ym�J����GO���._��Z�f&Fa�=�ϡ�����"}�X�a�)��]T(��[p���PHw�֏V#������	pY:<^)�k60c�8|�4��BU،Wg_��s�a�n�%���d?�UDhW�҉W���磴�I�Z^�sn�=�;�*��I��N-.�6O=ѾG�!L�$�I�Q
)��X� nhH.�a�Q�t-:�_���q��:��FIr�\�l���Y�ɍ�E!��0!���L�72r�U\�-�e�����'� �����+(~�	����v���>��1q�Ͽ>n	���a����&�{mڀ��e|��p��W��K��b��YC�N�'N���hX�.�=s��8yW��-#�P�t�R;e.6k�P�f�2�GX|�4�����R�F=8n��3.�<�>���Kxe�0,�?��v�N�&�އ ]���N<��ǠĘ��(Q3�J�LA�(Sn�LW�����~��ʭ��3ɮ4R�@�XϬu\�C��r��%��]�N��Ft��sa���"%)*�3�JDۃ�?;�,�>��g�dt����m��.nC����'~8z��=�ipI�5�Z*4�4���M|�?����Q*�15���i���<��'8a�Ll�jѼ�cl�ۃ�9f(���S����G���|ڈ{ߏc'^�u��m��6�_�����W���^���0�;������(d5/�5WL��{�iS�̇�a�Rȕ"\y�:��{�-A5"�J4\y���K�xv˚�Z��m�6��P��˔�Th,,ɧ.#�$)��)ZN2"߳��+��
nYVa:*��4��_�(xe2��]jhȗ����ݭ����t|�<�]<v�e��l��۱a����c�;o�h5v'5A�YB�¯���3u�ƈ�(T�5o����/l>`nLшJ��{�V5fp������BԼ	o, h�8���
�2`UZ=z����m�[�_��f.����ZD����W�=c:|�l�PҪ����3t�غ8�Bd�
Bt*7��\4Y�$�F`š$�J4�����.��G� jvg�3�f�r'K��L��<�"�4;+�)n��?�5<RY[��v7����5,]0��=NW���������Ġ	J�^&8�q(��P���?����,� �˴�NJ $,�z
�Z�����Z^�]#5|F/������k��B��b��.e���]�^N~����2uxF
MZ�T-�ЭC嵫�5}��r�8t����G&�$qR03u��Z(�5p� �\�ݨ��ƘGY	X�|BW��=�X�rv(�L&����Z��bq���L
㲶����cIӦăI����a,�n���Jsg5��R�� mZ������%N�a���m�7������?z֥��=>x�]j�J�P)V+ ��z�$��5$Q�y�� ����N6ZaR����
�/!��?�S�%�)Z��$�/�B��n�(�l=]*
��tRI]G�L�͗$�Ϧ�'w{��1E,C,Sig�Q�Z>|*7�z��H�$ϰ�h�[BZg>	P�N�B��������\�<ߚ�;�bi�x��}$������?��vJ������l�ǃ5zv�2��)�ѫ��)��B�h3�q[�1��ѳFL�����!1�x���u�,Q�T:��H���2�ZYk0����"�mnCJ�0*+v|��\��i��Ȯg I$���d��'�?G�ȫ�	��l�0�x
(D�{.��O�0� 6o���J>�˼Df3>0���h���|�L����K��tV�	D4��PG�v�4ĄuM[��wx�7�F	�
��l�K>���x��sQSi6�dh�Y脍b+�_1dԨ����;�Y�c�d�Q�[�j��6����6�%�i2I���>X���y�]J[�P���q:L�Z����BX)n)�n�˓��SKOk���؅GZ-�/c|�|/�&O�f������\ض	�+��<���m�ek�^��h������j���吧�x�>ue��}ʿ4]YT	�21�c���'^��_٭a�}�#g��<���x�3���5�a��C0c�.��.<�n����)W@d�ҭ�}urwuch�,�q�Γ��U�R�N����=Rv_=q�K�X�R�`,'�a��
����t�e��'�g�Zm|@��fg	� =m��c4���z7�C�b��7%���6e��R0p�$��SQX�+r�R˴�|^�x��7_q☑C_ޭa����3FM���6F���-jq����<{VTF�U���&|�H*a~�'�8�e,�[&�q,��-����8F�!-��	W�Q#���"��ƀ��7QCU��)i�/�I�
x�~�s:�*oD�zH���?�c�����<��3�ﬅNT�����P��7[�<hV�
Me�����Z\��E�b����|6/[8�ї���=�#?5e�/�j�"�a�mM��r�FP�4�ӷ�C�k@�cI^ �c�ſ��������?���RS��h�x$�Lx�\ghе3IV�Q�;D�h1&bw`�=�1M=8���֎���o�m��""����@I�3'#��.�� ���vu�c1<��lGr�b� ��ѱ��p�K���!{3�2�7�+	��BI�1b��-[8��=�RQ������d_�Ca�f?����x��@����m�k�3�J�.����s *��{��VW���{�L�N	������x_>V��P֫��G��ʆeo����R񝯖������\8Z�oy����,r0�&�RA�mNUʛ	��cP��=����8�(J%��f5M1�7W���Ο{��R	1�1�'Ti�&��r8b��Cy�����,���*!P�,F�W@my^�c-�=��0�+��R�mj،��M�&O^e���a5�C��5S�'�T�?�\d�U(�K0���،�/���D)�/�����|�7^!�iIN�XLOb���n X{�� �I �A/lDgm+�����=������ҵ��0�/b�[����,�vVD�c����������{$��'ޗ�O�>Co��ϡ0m��C'�u�-�j���0���%m���w[C؆#WV��8�d�E�]dc՝�p���ثc��^� L�����T�|�t���2�F��'(c�c�<b��8z�5�g����!й�A�+&�1��b	l��3)W�򐽗�߈��F<s�L���Km���`��X����`R,�*���롇��F���;>r:�:�ރ�/�OY���%�jh1��;X�%��b���F������=��Q��������0BW��$�e�ni�q�=w"�u�W#h�{7P\>b�T4��Wk�P�� �7�6u���:�z!o�IBC҈S��\5��H|�Y�Ӵ�����0d�	�]���ų0n��8f`/^I��P�X8w>V����D�����a�3X�a�~ElT�qg�!L�@�h^�}\~��i'��0*�mhp�f[ҍ�i���7���5����a��I�֩C�W�E%��KF�P�9�N�����u���p264E�b��8b̵�W퍂Q�*$��\��R�������q��&���M!�`v�C�h3�_2cƟ�c�F�g#O���ebѼ�X��[r�bt����܇|DF�N 5���GLG�����`i���=��%܄�w��0dEqʜ'��1�&�0D��E���T�(,�3];w��^K��p���O��N���=dȉ�B	�����3�.�c���Y�����z�l�1�I�]�<ŗ5A���v�n����DegK(�d7�&�ml����7b�*���T��[��v��y�Gv%����2��l��X��s���1i���dInO���<�J����U���ѹs�j���	�K1BF{^C�R�95e��,��]�|�^(Y�`�Q��	A`�K*1-���~��8W%���zzVP����%31n�98f`_�0�"<±M,�{V�Z�89��'�{�=��c؈��}����,�P2
s���u�s(I<F�c�}}k���h�a��C	�1�4��蓙kT>���Fa�܉�Թ{�����/�a�㹫��x���t��]�u��rfM^��hJ��	�gF�d��c:"����� {Z��C�a�2�����lØ0�,;��pl�*��[�Pr�\�JA[ƞ��#>$a���
�_(�q=�8�������+���y���2rҼ?��0T��鞮sa9�,K)"������F`��ɨ��M<���ɰ)�#GUB	�4�{����O��KGHKPTL>s�O^�c/��l/�*��M�����KbY	��'&�_�0,;�\-;(���9�_<��� ��%M)��0eo���j�W�{��|.��JP��a#����ֆa��v{�6Ɗ�;y���j�a�a�^=�1T��:�1�\��2̝;]:u�K�{��#b�h�+WUɨxs��Æf�'-��/��L/A��&��$S@B$�e�QC��;��v�-ư��w� H�)2�j�~�B��w��/����$��m,�V�z'|U�=��r5f
����/��.إa�Y��QUI�p3V�qyn���C�8D��G�9b�ܧ�b��P���Y$WFd6�mF��1��l:�q:�Lnd���0��F��tT<���Y'�de�7��s�i8��d�@� �|��}L��z�8��ӽШU#G!�te�k�#LH�T�S�J8�a�T6���vu}��q'�9���L&��،��zl�3fa��q��_���EQ9�O�馛��悔ޝR(����~�1�8�7l�5t�$t?�:�z&FW*��8�!��k���RU$��p�%��vø���O9yޟ�j:�N@.��%�!�/n��gxeŵ����9EN�"L8p�Uh�7�?<�1Zݡ�^E�E�
A�AK�n��à��(,���	��&V��o8�G���(�(h\Z,�{5z�$�P���k��P�ʎ��ŋ)#QH+5ZQ�$��8�r#:�#8�6�����e@o�ۧ^PhZ��]�^�����o���JV~�μ&O�����=G �+W(��?��ngM��� ��p]�7$���{�kk�1�m���؉�L�����$� �M�8V��	�x��o��A�l����2'�B(�Co}:c�
�o�M��\����gJ��􀓿-]��⺃	�
ƺj�1QT����I�P#���![�c���H`}
�����l՛aI �Qqh�z�    IDAT���_��@�d�-\�����m~�GT���.D�Yu�Bz[��T[ �:�u��0k���|$�&���0�$�4/_4��=��v���q@�d�+`��}#ȣC*@��`��HBƜ���t��bHJevo�sۊM���Bj��mo���Dx�03Uȗ�l��I�0��I�������A'���+��Z��L�� /@п��U�CgF���/�1#�V�^!}�+P��x�3�*q�2�
~��c�^��A��Q$a��g	L��6�hv&n��}XE+�Ð�Wo"M�,�f���<�F"x��͟�,�ui�E)��ga!�D���#��,7�\��!�/�LjP�CGI))<]�O!?�0��&1 ������)gU���9�{镴r+���*A�:4M�\�҈i�g�[H�j�c|��j�ؾ��g�,����6?=!#W��Ie�FI<I��\i�q�;k�|��}��F�rAC�)� Nt�Q#Ur,ͤ��y��l��(��%7���![�fkP���?K�6�} �t�pG���2'�݌�܎������??	I�)����"�|aK�Q��G�c;!�8A�DȈ6;�b�x���R�>����+8"��{��q+v����x�$4
�z�X��uJm�6@������0ڄ�jWUR1{Ob�Z�Qw��{&�+�2d�c��I���Q.Tx���(V�� ?R	�Z�yTF�����.�X�����_p����l|4��7�#Ij�O;i�I�T1�ib�\�?5*{�X��%����0	K���(r΂iā��(�[b;3�؃%�n4.A��Z��\v�lE�m0�ۨ0���+�xbl�c(�yk��&�h_�+nq��i��#n)#����f�Ҫ%��!��̡x�=�:�L�S����Gy �V�^*���X̋k%��l�k�ZO��c=*wGMg����Crbe�!�8�I�+�Y�0i�'����sɼDȢ��Ğ�>1lz	~�xO��U��k�O�?!k���%��Da ^)`4y��z��%$w��hLP�x����7Oo�-q��J�t�+Hnl�	�I����O�ѿH-�<�J�8�����[��s���-�S~�1���l9^Ib���mx���-�ɱXFȄQ���v9ȚG쩨%ƽ?R�
���q�{'�xw�bj�4}al��"U����h|��]�֯����cH����ю骂ޫ�͆��bɆ$�'#n�8����$i����\kI�*�H������_�Ժ�3$V�5�0�¸�&�^�k8DV��	h4�c�v%�xr���Q8��p�̟a�+y�R��^J����7Y�ja:n�����!���M����r��GM�G|�$�k���oF{��u�j��Ee�-E� �zc���B0�`�Eۑ}ng�۟���M$y�� �a�?B���a�aҕ���G��� �Cl��&qd퉇��J��1q��i��ai�����~\�R�Dr8Z_�T9�G%{}�o��j �S���{�>Lؾ%�r��x�v ��tQ����j�I=%� C69 |H���sw������#_�8f2]�ױBH�[�Z�&�=.��	��!���7��"Yud���?�*�/���]hh�5�RQ8�T*\1�������D�5)��sԿT�Ί-��Q��ѹ�����i���%� Kj�4��%=^DR��� �Klb:�|���x�<I�J�h�{��H�2C��[��S1h��e�P��k@]M��7�(l�WjĖmM��J�lMg�k:	�g!�����0"�?[]]YH�]=$Uٴb⑊C}�@�Z!�X�������
ٶ}v����[�ў����D�/u3x
�z��E���!���FO�|�r��b-yF[�dL/�=���Q���lpe�r��|Ԛ6�}�W>|���V:=�b���PW��|�lY��"��s �p:����EIKAKנ�(p�>�5�@k�QM҇V}�=>�V_�ŃQ����`_��a���}G���2��˜C@0��|+�B�$S��M0��	>���J�RNO뤬-��g�B�LF#iH��뜩�ѻS5>~�oX� o�N�C�9��?2�(����T��o���<�L�|*`T��w�G�����ed����2wQ��˅�(UM���V���*��dUA	ͨ܄��%�b�P@�<�����ٴ��5�$g��)�+w�U����ln�)UwT>/G��IC�|�q���m�z
��ADb��ql�?��*-,�n8�����r�=��A/�?������Ko��OEV��hI`��#n�y�o��\���y	g�v.��0q��[���g`ejĚ*�q�h��jy�Ʉ6A�WtYHRO]��=(
�?�+Ir��*+I�e�̕�Lg�/���wa)�9�P�V���/.��'P���z�s�L�, �ƢIĮ���� r|R�U���^�f�\�V�JbFd�7�ؖN0INI*�5�%��n	�TVi#��>���/�A�{��A�^��|�����8J*���x�u��w�Mx��_��3�g�ES�F٠�ԅz�Xצ��LZh��*7��L̻U���DtԷ�[��͊m�u� s��?�.S�(f ������Yp�(e�~��$6%gUj��G�l��앴u���7Q��B�D����	�1�����q�_�~{w�
#Ij �8VUa�B|�������Kg!_u0rf�����_�� w�L�M9!ZT�_:��D���t�6���3p�����?�S@A�n
��KQ�����c��]�#�&��Il�\ ���ab������p�����썜Ü�BT,�4�� i���B"q&$ơ2 �2��HS��o~���z��z1��W�荰�֌4��`�y����t���+f.�~ρֽ?"�k�1H�Cq������q�=YjnSK�=9F�㎉X2
:v�(�x�iȌ�;���ΤMB��0k�|{��(��-A*��ܹaȅ�E<�� �����b���~�c�d�_.��tQ�	��U|�e�Ðe|�ylj`�S ��H�	�-Ǐ��)�6��}�L�N�)���mt��*aAP��(��sE�.�QS��m�]3V��!Io��~G+,�y��T-�����a�x����w�1Sh����v���6�q���׈I�~�6�N�<�mKf�W�[#5�	���J薘`q&@��isp�%W��?Mz�"\߅ǐ��������۫�����_݃O��A�=�8,�,�>R�'�$7R{a��#�SÓ�2��m�p��9_�*{�t.���vE�PVd�%�?(+��D4QRV���e;C�� j^��<��*��x!�8pX~$�y�XK�Ca�:���F��}4W<Fblʩ�u`��6������NB�q9	�j9s��@o��L-�{
���l�b��K���>�2Y�yD����qV�9���c8���Qs�D��hLt�<aq���0�fv�K�{%1U(O������б8�F�kz��;�H�J�TX�e)Q)x�,qE�<�����̒i�l�0֯�0�����.���Tʉ
�����𑳰߰���u���a���ѦPr�̾n��o?�I��� U�lI,�t���\u�m8���1�r��̮B	2��rR6B7��Q�������{�ۯ/�(�u\��\�����4�*M6��(�"Xr��u��1@fç܀��y�8l���,n�U��T�Y�HJ,)�w�Ie��ft
?�P2��0�O��&��S���)�:m[�����=�&�z�TӐ�_B �r�Ģ��S�Ю�+7�[�ᔓ���C����7Pg����&+_x���	��`l�2�T��0X	��rK�2<8����W���'7@��,�=ߓ0��_@�i��f�3[��q�R�_�#���z���[ߌ��"��Z��\K��e�Qs�Ua��a$ɧ��Y6P���Uۀ�,��C�; ]�j,E�O�!S]+B����1��_��E���F1Jn����F���Sy�Sǎ� �5-�(���i��
��f�N9Jw�c����CGLG�n����W%1�"˴z� �ӗ����!,}("�"qMv?�u��P�Jܔ�&Y�.RQE [�Im�F.q�X����<#�����G��'�1�J�T�'�妆p�;�p�1����UF\�)Ɩ7��7b��a���0�PE�43�|��!o�*��e4�������a�=PH�:@�!�_���ʫ�[�y��)�^[^v����&iZ��%�T��(Wc�3;�Aя�1چ�K�`@]�~��iP`�/5�Pq]�S�'��G�N����W�Jꪥ靌��G���[~���?���3�e���mT������d+�&&9Cd�&����ܭ�����!����o������,2��`��iZ	f���9Wi��%9��~��_�EU�e�%mB��}��?9i�Ͽªą�N����j�ap4E"�,t��`�/�䳇�ic+({�M���b�Hش8�-���dd�IL�֪z\T�4��o��������a�ᆊ[���2�ފ"�H�iőE�7	��7�9�R��V�4�?j�a�kS����14H�[p}�:d�?�'?�+������:eɾ�<IO�j�f���_�lF,�IB��k$i\k��˯��y�>�n|�Պx�n�BtO��+ K����&�G�v�fcG����X��4[�ߘ=���\�����E�2np%-��z���rو�^m}nw���� ��Ð:ݴ��`�l��>O,�	�;���I
�x��vx�U٨"_M��yղt˸[��Tǵ2���~��50�3�^�Ԑ"�Ꮠ@6�uGu8��jng��Ƕ�"Z��a��0�bzU�#+�j�P�/iKc��+��#3���=r���s�
C���l˫�D+�|H1�[�����n���Gc���W9��1�V=�u�\W�h�]��n
��P�\��X��/}�����C���Iw�!�C؄�%/��NƆ�ȑ�Q����+���!�ǿ��[����a4-[8��ї\��<�#珘4����0��Z�.�d�2����F��a������.?�/=Oe�0 �yp�G��8�`I��ۣW�mC��r�/n�Wf+��x
�?gMX��A��+�r���sD�p�:�Q&�9CSp�v��4�� �M#w����WV��/��6z���7O�Ƙ��ڭa�}����<�_�aD�ZG��-�v�����f6��o���ϱ�+`�]�d�Z&�n<�2)�^��*Q�&NB���H]���O��VǼ�Kqǯ^�ާO�'�j����/_����<M�`�(i��cH�о䳨A{0fh���?k�>z��)s~�V��4X���p^)�
�9E�����1�����ֽ{�Mm��}MҢnG��&Q�t��X
l�� ƥa8�٩m�H��6����Ŧ��Dyh��R�D=t[2���QU�s[r�{�8U�+��@��媅����A��4����C�Ƚ��%�S�*Q�A����
�����'x��Yx����l{�9=&�� �l��{k���Dmߣd���웴�iKF��n5lT�w�s(���헷�c����ᣦ̽�m�����M6V��i�BP�����;�G������o��x$wi$��ÃκL��>e���,9�⍕�t�yʓ�G���-˔�J+�����r5~�ԣ�α��� K�jx&s3�+Q	�a�Vj�$��S���;��:<Ɋ�����}�ހ��	������ݐ��M�jn���H��՚QW��,����z'5Pn�TO\�;J4��ka��n֜}���5U�W�}�7�]8]eK\�z���a�(�勧}�ҋ/X��P���#'Ϲ�-�����DÐ-3f|&4K�Ϸ��Ƨk^�|�����X��r��ϛ�a�Ð�;��Q�Tqf	�o� ���v�� Ҝ��O�W��7?^�,��5ٕ����H�u��Đ��7������rr{&I�QW/�}\���s���Ƀ$S���-�TrT���
!��(7�R�6t�>�SKf⅗�/��Z�Y��0"2*aek��{��Y3Q���C�J�b��!�S1S������\y����ڔc��0����`�.�*ӸBHè-|�ՋG���b٪�z�soCS�Y�q�z���o�3�^,au��Qml�y��t�Xh{����T,9Q��]�J���t²ZLՠ�i+:�BT����f�/�_�G�2KpP�c�	���G�1z����W	�����Z���ۊ~}���.�N��2��9��ٚ� �S�D�V�!�C3`�[ѱ�!^�g6�!��5a�|�x+np��#�$�d_�P���OB�3f���a���V���=ޤ(�O�Z��T���e"DI'B]�#��e�؈����B�Th�a���������/���� l
�����ceR�Ls�!��-"]���et��	����Q~�Y������j��: 5CH>Bq�
dGa˓W�*�/D�� �H�N�JRړ�=����3�l	2��!j�D��8�op��*�@���FM��ن?�t9�"˸(�}|��L
�|c�Ks���g�B�ϑ�.׸-�V&x��R�hO���,���2s�'+/����:�Z<�&����K��,)S��GU��l��Tl��<�F~��#�ڧd.�1NL���������SK�3���F���c8吽���"<Q�Z��
����Pf!RnqoCT�X��/gl'{ �����w����q�������1&�b(~�,��Pq~{sk
gz>JhTkE�4���V\�	��1��E� ꔃP#q��b���Y��9��Q�x��Ͽ�^�Ǥ�VL�~�b�I�<�%�����^à��*�(q���,���닆a�3q�atw6��Z&.�[�a)/�O�Ic�W_��OE��`4���g�aPK��t��R���Mq�|3�j��{y����?�+w/�/<�/���g>{�Vӱ$�y���J
 j���Kzs�҇0�y8f�upS]QD5�	�m	�!ق�y��D����Q�����fb���qD��Đ�+���(K�Ͳ8�[:硗LG���
�g  XՈ���0V��M��6b�ڒ|��ÈҒ ꑇN�:���"\5c����2�l8i�\�@ΦӢqFؘ�0sҍ8l��(���?%�Z��� �� S-g�<�n�kR+,*��N	G��1���Y��[��G���	�(R*�H�cW[����\5����W�u`ظk���?ǠS`v�m��HO�H|��4�H�����������:� Kⅻ����g��=��q�� _R6:�Ӗ
9X)�G�Dߋo��c |�D0�����	o�R��*�l�a�ݎ>���TʄdV4hiA*Q��s�+]�i���!��E��B l8���{�42Ӭ����+P�P�b>c�Sº��wPnB~u[})�z&�&��CD�Y�&X����ۯ��?�í+c���@$��ċ(�:�PP���~Ç�:��#�Uݱ>�ê� b}��x�����"nC�e��<^h80�[�����2�ǜ�c�)�O��f�N5B.NŬB4,'e���	�N���X�kx�����H��ٽa�Rs�]f���!Z�:��8�'U��y#q�vXF'�_<
�ǝ���<����OJfˠ�L!W��W56t�C�,�����[���V�|4�q�3�D&�Ze�N�@JREt�����+����2#'\��:�uA�\[��:��/���}�u\q�B`�����#N��&_�Nu�rQ���0����h��C�dJ������e�L��1p?�,�Ejy?R���pH�����G�B��C�1PV�Rg�$�D�uC�-I��-����&�Xq�CGM��`[BI��j�ֆ�	ʨ�c��1�t��8f� ��BK�p��zI���L����s�V�~��<|��}���ʴl�'$�����Q��/���c��*��	��6`�'�b���QX������_��i+���y�>�Px8�>��C���5hU��T�@L�    IDATv��/j[�|YÐ�'ӗR�ݍx�q���#���n�t��?�I�R�%�w���Y���л��KY5v�cm�|2�n��ضy�{�o�-�6@e��j��*܌�n�p�@�Iy5�F��җ�q�&���b�������y�NZ����M�v�N���d�@�i1ތ�����(5"��r���I+�a�6��W*ɺa�_
������ �,�"85]��)4�
"����YxLwiINQ�!�6�e��uQ���f���f��yU��'���
b��oy�3�j��+<�I�#�DS�uh�-ø����9y��m�I#�$�$�gV�#P��6j-]䤂����#���k:�.қ����0�ڽ��7kD��8M���1��*E�|~���.I�uN�q5���eW���Dl*�(-�2[�wcU�2�l;KXI�H�6f*��\�L鴃b!�T�VDg�b�Ȏ4K�)x�D�7 y�������G��v^A���0SҊ�����Q���l����Ɗ͒����7���8a�x��?z�Isi�aHqse�9�/]I��V/�aK�wQv}�p�TZ��n�Uf��e����7��s)�M^�@�	U+\���0ĿDj��xϗ)-x�Z�a�@x�Iƚ�����2%"|#�J�*��jh*9qY�����%�({�+.SC(�)�B"��i������^]�2T�`"���҆�D_����0�4%�,J�}��P����/H��F������E��l���\*�o\�p�=�1����Dn`+* �x%�)���[�JV��(���I-#�c�z�W-%��7�+aS�J@��@�`�l�/��YJ\���c�8�Ed�iY�XM�1����lPF�hq]�G7
�!��s�َ��[P�'�<d3�_c��-��n�3��=��T]VAɲ��	˟���YK6��G(�x��j�RN��H��*�P��(��0V���٣��{�����"�3,)����Q��R�,d�Q�U�M+Q+Hq	�j�t�|p�4t�!�����K�-���*�)T�.%���ϝ<��|��z�ghJc]QI2�(�6��&�@,+��Mtۅ��W'7�"6a�)�*'o����s�PQ����w��~.{8�c�ՠt�(OxL���*I���>��-9���B��)U򲖮g�c��0��<��6 uڮ�|�����yLɖᯠ<]�Cn %���{�*�bY����IOD*'5�J����I�9�O���I
���~�����8�I�TU�A�'��.zn����JA��Ϲ���8�5uSI>p_�]NI�ZA�c2:E���U6��A��[11q'��/:|�ra��Y�}YT���vF	;�dُ�eΐ�0�ސLSe�[�S�>�T�J�/���=��ۃ.��$TJ�"P8Q-���"5�u2�(�p]��Д˫�C�k��#�
!��Qln�ϕ8 �R���U�r�I}c)���u't��l�5!���GVg�Z:V�_DZK����;#W�s�0*
קw��`%
�+wI�It�p�M��JjE'�	p�����P��KlYS�_��JO�PjY�đ!��,�[U�7׀�AI1Ű^P�l��Q��N#�z�����qJ���W|��A�("��bI�%���dm���TTjB�Y��aC`��pR5ꁺEX��M�$E������VXB�a�{�Fs���	���<)���q_Z��Q�b�,-M��*�JY�dYF^N��ٍ�A�.��r	�Cɍ&ľ��d�#>������_B�LŇC-.�������+�oǥ� ��j���-t���lM5�%5��$��D�v)�3�BP'�7cl+�<�n I�%�r�H��������D�c!�J�c��X� D���*�8��\��ݺ�Cڑ!N�4:o�/b��*E�y(�s�i*GH�����|^Z	ZA<�DV+N�K�	�S\��+�2]�d��=w�l��x^#,ǂg����&�i��\��|N
�b���t�A)�jH-V�|G�%a��'�����Z:h��fb(���$r6+��0@���s#hl����,XF���Q���"��(A�oy���k{��C��*}S��ɤ��,&�erZ;B���6C3#)b"�M9�BH�g�34�]��r*�R2m��!� ��u�䉬�,j���؉T@6A.�T��G(����t��ư#zL�y�"�� n䢙���� �T-rVHY)��y���#��p�ɕD����p�+8_ �+�'*[�Ԭ1|��,Sl'R<;L��������\��Y(�Bx�S�\�衐;��P,Y����0ڷp�2k�!koE���L`*3-�F�F9����7���	U�#d�.̭nIT!&#���pɱ)�<ܮʺi�2Bu�٢���"���	�R)�~lp	P,�^��Z�\>&�
q����p#���b�ơ�eSY���c��)4E1�t�B�P��R7�Ur��*�&هm[s�4�L#Dѣa8r8��Ӏjzٲ���PE"�#�@���K�BB}i�E�?�&���P�&�ؕ�X�p�W��P7 ���F������&��0��'aӨ��oF��	���i�:��YzU��CN�#t���e��\C���
��ѳX�M�Ig�d��r&2`���.�ha��e갵"
�m��nظU��u���T�[���5Ǉ����a�a���(����1�����Q<�L�Z���zҠl�% a�C�ə�B�sa��<�xՖ���|��W�P(QۡNr(�����\tѣ�^H�r��l]�X[_�2����پ���|*:B���b�Qx"��͓��B�ۄ���ǡ�Bm�Z�������+��ߗ��G(4n·���y��?�U.oP3��zϬ^O�@��p��4��طe�ې��r���W=�[��;��ף�Cg�|�x�w�A��M]R.z�쁗�[����c�늌��J���{���O�0�����*ui�������L�]Y���]�RN�����s͠���c��zⵕ���ǀ��q��A��^��	��� �WF��0��1x`?4or��k�fK[K��/ۣ�ve(��1M;i��h흮�
��*�4�f��_@��Ƀ:�_o�<�V�
|��s��n�� �Y�a�]t�i�k�:|��'0�4�[?��}7\�����!���%Nxc}�B�湗�i<�*�IT�KRjVa�bȡ}1qTo��%��Qk��o�����⋿���	=�6�TzX{�!�p�/q�Q�b�y=�֫e��� �����;؝��h0P�\��ȕ!"jϬ��pr������G3�E��
Qӧ9�����{�O1�GCq�`/�=Ė���l�r˳���p���!p��/oA���e���^�V"����Si�k�1�i��3NڳRs;�:I��ت�Oվ�����}�&e"�o�ms��+n~~�%�Aˮ=/<�1~���y�yx�X��x�ݷ�ǣ�OŲe/���`�Kw����7�?��&�u�,�Q�A�.�uK03���������O���4�P�fk��z�zv��o�}�æ='?�� �&���&�C���ptg�x����p�����b՛y���ߠ��P�!ym���zbA�"M덫���s0e΋�|�m�+��߽Z��F��� ��|�࡬G��s����Q_���?���A)@�J�>[�T�!�7c��Y�}�y�hm[;@Lڃ��a�a(JQ<>����5�,7c`�z\x� �h��t�B���ۀ)�5�t0k�Op弋���>��~�Щ�߼?�w��7�ޔHےK��-f��t�s�˿�՛�j$��������]0��>�A�k?l+z�ׄ*�N�����o��Go�����ƕW��{�1v�i�h�8��#q�{bܔ���v(P��C��o���������0�(����t���Ȕ�a��`d��Kđ}�a⸓1z�C8��� �ࣿz
MZ/�4�L��'��ϋ��{��#��R���Y�w����� U�EDε�+��b���G��`����� <����۶YI���Y�ڔJ�*�GCC�p�)��ē:�򫟄�aXv=����N�|����Y+p�Q��ck�v�68���#�����^�S�d4~��!X�6��~�
�N7ԊDX���Ȱ
�n�)͍ͮ�p�1�����p�#(:�6�[ؿ�<_�z�s8x�!��I��}�r�y�x���b��0tԷ1�ʟ�SO��'�b�5� �=K����8��#pѕ�0LQ8����4�SZAHIM�oވ>=:b¨��r�
�6T&���ߏ��Fc��?}���3�����em �~7�$̜r/>3{!��yW��,Æ�!#����c4ߵ`�ɗ���n=���>r��)s�i�a(�E����I����3~	��	��Maܘ�8��G����M�*�0컇�G�,��	L��,<�Л����ix�mx`��~��V��-�p�����5�g/�OwGFKJ2͊��`�-s��T��{�`�E=1}��0;tG��ѷC��c��ᓟD���q�=qͬп�>�1���ﮧp�ȓ1lگ��O��N��u7��:[7�ǹ������a3�v_�Q;�Twdc�8� ��G@=ִ-�qż�q�-´I�`�m�����̪�Z����93��PFA�!16�r��(j�I~#�Ad�� )6�WQA�A��$�2 خb	2���9gN��f�ooa�k�y<O���o�o���U�������ˮ�h�_��폂�C���hށUs/������� ,�#P�H"Ef�^R�j��|�;��,
=4�_'�|��lF5��&^��lĶ5�u�ނYS���;_⩗_�-�]���X���֡.�桤���؉��(�ɜ1���h㞧6�t�f��D�T�7�@�9b*sp߄JQ����s���*6�F$�Y�%[8nZ��8	���7O{��è���
\��Ӟƙ��E��;`���?�d465`�X���Wo�)d���Ty�H����$R�Ԝ<�&����8��/ ��|��qr�1�:|!�pg$lb!���fa�Ⱦ��ۘ��i4
:uA}���i����w�+Y5��T���dT&$;I�q��ۋ/����w�植�N��l��]9�3z�聑����{@m��~��x�=��e/B���j�6�\$����/C	���5@���WS�:�.+M�.��^��/���kZ�9�ǅ��":�U�:�L��7���=�`~'��v���D�;�9�~֯q]���C aǝl�R�c �,����&�M�g�'�OC�)1�@N�[��_����_�� ���8n�Gu������/�@���]w\�ʝ��-@^PCYɚ��G,�h[��A�h�b������?���x�<J��F�����>5�t&o7�P,��%e"VW�ӎ;'��S�s�lM��w߆�`j9��4qF��(������a��g~->(V
�W���슛H��P:�+�Ӊ��M=I�yU�����il7"!�\t�! Yc`��j|�����'�_|�vN�]���rQTt$_�ݏ��~�Aꯨ>���d{�
�
EE��A�� %>oBN���\��t����2�G�>��O?a�?I�L�`%�����X��Zl���d�p'��D��g$-��u[�O�.֌PN������V��c��C�0���=sU)Ȑ�=��a#�#��S7�7Z�P��H.o����Ò0R-h'�nG�D
��|dH�D�3
�$d��*�����,�]e���P�ށi���g"9~�$�k�!H��$� O�Y��h���:k2�0-)�x��.|2R��P��Ɍ�K�$�3$�C�ɢHc�g/�t$`D���#�!��`�a�`F"[63�8`��z:Ú(�t>Ӏ�hJ�hױ�Ob-[��Z\͖���,�WXۢ��j@E'������I,����S�1�%f�4$�..�O� KBʰ�H�Y��:dL��.)YZ������=A�I��_h����Q$�Is�n�M���1H���a�SU0�Լ�?�d�ivj�z���_VGtU�\�J8Sj�;
�J�+����룣��b�ϝ���$��}�D"P�xV�	^�t�NӤ_J�K�=�ᙓ.1��~��č��L�#E�J�%�_P\�I�E�uN�3`mr�9V��S��G �hD�~^i�����iK�(E\�J|�t��n=��A�Fe�!�q�Rw�J1D�#{�l�4���N��7��*�ihhDT5� �GR�<$�s�1�p�Ej��bP��$b!��4!�#��ޑ���Sy�&��V~��AR��X:}!�u/DP�{���1�5����o����͒2T��Fm!��4L�:�&�i@*�+t)H1UN	�)�����P;:'Ľ��� �cW4fd�dd.���E�r���
� ���A��X�6��,�6Gy"�VEgԃ�y�Ds-l"f�izNw(�����<�"��$�!��7�0�X���Cد ������)��Mք���@���}P5���BGSFB�{o4e迉��f|��+p��/�q�o���q@�X�xŐ!��~��u���<ڣ&b>K�M�r�B�I2����&Rk�L�KuDVO%qŁx�|�D���PvҁBH�KLx�� ���[f�F�IO h5��s�t����"<j6����oݠ
�C9��~�<xD�<��A����뽨�	(��P�l&Q�y=��z�A�
�����T>�z<*)�O�r��i� �
���#1�I�>��4�KV-wׂ���]�8��/�:�;_Bp>��f`��AX����hx���EZɛ�"�[�E��ۣ- a;�G���+��I�?�I�a,���&�@��rX|:�:7㍹� f=��`n$�H�o����Ť��Fd@m��Jq�)��QKF�ʢ-�w�s/n�!�(��D�R��jT���J���Sg<�rIz󎞡��AHw�^�g#�+�e��&�q?�W�+1֔��E�7�c2��G�n�@a�
}t�/q7L����B��F����z�|�r��@��:�o*���/�Y��v�/�NG��)���v�N��=Q:�UR�%oefP�Ϡ�ڃWg�dvv�}#�-qc9�<�n��K�N���'��[�#����x��;Pc�:͊
_��M/a�ߖ��i1��j���9�����<�j�1�aĔ#��d��1�Ɣ�]�{&_rݐ���1���l�]��j�=����G
���$��AnN�H"�I�����������V�G�hE�\(�&�i�Y�G��Q����
ӟ� w���Q��4m/e�\��#�nDAf'�?8�l����+�-"F➠6W���Px�(��	;��,(�R>z?ϣ��qB5bϣ��ֲ槫Q�z)T���\2��E�m�SN��~���Dq�	�OX�z���l/�^�Ѳ`��K�J��,��~脻l�a����]���*d��i�J�Sȓh��2v�0�ټW}�{@"#�%T���$��΁T����v3)�������8��(�[[!��2��jtqvc��I�̯�'Jw[���d�Fb2J)�.��ec��� ��c8v�M�����yXWI��9zқ����j�3��l�db�Q�~�M�DW���^�}&,D����L<�����y3'^:|蠊{�%+F�������`��#���?�\�d�t�eu�[
|��1����^5���9��AWE"o4�A�:�R�T\� }�Z7�=�nԨG0��x�i @d#���$�G�N9v3
t"Z���=q`� �m��N]q^RC��G���Ǣ�	�!-�p�U���*Hd��<B�6ȨLGF;�{�il_�?P�Z��G
�b���)
t+-T=�b6�|��a1���,���<y��g�gM�lXt�ڃ��c���y�bh�����2���
6��Q����C�l��b�s  �IDATFِͪL�9̫�O����nGn��ۓ,��	c���+� �H�=�N�)G I�*�]�(���3]�`q�a�|,-C3�_a��ɀ���d .}��%�qR��ИHs
H���=��-_����j'^6��)9����<N�x�]�tw�����齿b��_Q��4���i��B$'i��k�][��̀e�^��L-DѠv�ek<}�*���0��gM��"�砆�p��qC��5���Ὕ�C�C�TB^sg��BQ������nA��5�[u/?�{��*�s=��B�"���9���$ʮ��
���l}�ށ:�I9��*�àݤ�M��J�Ŵ����x�̀�`6{�7L�������$��h2&���;����|��)9���^,A�S����a����"D�8��]�]/-㬈��4HE5��KW�b[&��(�q�5�����7,F��6Iw1-D[�.?Ʒ�h�y3�\6|h�k���ax4C%Z1u�N��o.it�g Ό�ͯ�n�}�Y�����N3f݋�Y��F���rc3�=J:����W;!)繴��+ܹ P�u\�#�k�l��x�-�U��l�d�c&��/N�	���-U������/�~�0.����EF��`(٘���<��l1F.ZP��*�~���HN��^��=�P(���pn��FL�2ŕ�d J�:i�#�X2$��ګ�������ߑ���c<�h�ء����m��
�8�:/t��n�+��v`�Q��g��(<:T����.��nhsH'���Q7s f_�d��^툤�+��jyj͕�o����i �đkVc��[������N�8}N;����"5�n��TTn�r5MX����@���c�:�^AM̮�0���[B�(Ix�����a5p�̌�2p����ɇ����ݜ60��1"���.��	}&>�_� 4��<]�	��e�fN���磋W�:����b��9=e�m�l�@P���IL����"���M�~�Hv�p�6�{/��LI�SX�2"8��<u��q��Q鈔,x@|^̊~���M��l�#Ϩ��{ou=F���ɓ�3�N�͚�A�f�uL��fl۾�5�L�.���aPZ*�ἴA���D�{A���%a�?�]lM�㟞t��#77Eg���`��񮖊�j��c,A��H7@���U~ �.�X0{��MW�Y	Sr�H��/	������p����QQ0i h��a�z�(N����F����E^$��:{i�h���PF�낳�ގ�0Zȭ�}o*g*��pD~b�a4�Q��>2�� US1f�H�:�'�3ҀM�O�6_T��j!
.��ǟ���m��6E�Dɉ����.�,�� d�a���M��B�F����9�AD�~�-��il�1��[�j��`��`*]�{�c�����h�oo�2��0�g�E-p-\�l��3�5�Ԡ��y>x��H}�(��"���3j����>�OйK�)��2"]ݼ;V- �Q��������Da~G��I9��Dݣ��Z�;�N��af����
���^����yX'��݌\���a�vL�q��ĉpꩽВLs5����4m**+w����^� �/��O�+uk!��%�'�*hH��->Z�J1�~�<����0��н�C��8�&��Q݀&L� �|u���LZ�G	���[ܶT�@G��3'�f��A�������1d���:f1��B� �"[%4�jc�H)�$2v�8���EB��x�ILA�C��+��o+�[#���m��~��ܾ��& J�R!?JXr����Q� f��#�[�`��k`�<ͮ�1����(YM�:��D�8F7�pN<�R���ɓ��˯��Ћ!��oJP���#��ʫ�z�5�����a!�ɼ~��_���|���WCs��~����׎'ۉ�1na܈�P�[���,��g�{�Z$-���j*�-�د�x`L˼{n�p��?���hђ��f�;u�b�!�!���t�N.�D��# 9̚Gmwj_s���W��p4��+��ހʏ6��:���D�@e�4f�1y9y��Q	9e��~�.|qT.k@�N�f4�"X�|����KɃ�^��8��g0:-��[K�si�L#�"��O�N�{�Yl7�<���?�v�r�(:�/�\�L�EMTQy���� 4�]i�(�L7 d7a���hx�9 ���W��W%̝>EyH;Ҏ��Ҙ~�T&���A��:f�+��˹/��5r'�����W��X��RR!`G�<<��~#�^u`������J��=��腨��9�XA�H�
zE	zBUO:k�<%w)PGn���72�US'����4�15ۑ�݁�_�q�m��|�C3|Mq�hV0�ɷ�)
����t?�$�I��a6\qxyi���T�aI�B��V-��ћ�h�4�4An�`����[;���)��ၥϠNꈌ�"��1m���w�*h+A8�#�bQ<INQ^�c#�qXB��d�64�4+�;*�D�ބ���F��iX�j�<,{�%Ȏ���g\
�[�~hQ0����b�i�6\�+y^nⲼ7Q-Ւa$�Ϟ��`����2��G��^�Z�0�����|��xR\�	�G�ܗ�Ӄ!"[p�A@��Y�rXݝ���P�8|�ǥ�uC'gBH!c+h��o6�l,[� �a�*�Ĕ�� �i*�*n��%ua�rFES�=̀^�j��'�x��_��_DpT ���3о+V��5��Ѣ��&+H�M�ׂ|}2�Z�Ȫ���b�7��N�L`!��Q��Lq�T�z9?B�j�?%cd$ah��Fg��h't҅�#�|4�R�\�LT��V��X[>�c�wЁ�K�K���Xt�臱G��L9��vQ�d��K`[����e9�V�!PR:쾴9DWd��Aq�����?V����n�nD�҆�X�h�Y_��Dn�%aD�C�0!�e'Y��[{o�%u!yo��\U�M#�To���A�b@�؃�����SKӬp"�k>m�6�H4�aPe�1�d�Z-n|�``�;:Fż,W��`��~��A<]�%�"�AH#nA�@?Y�Z\�S]�j` !��Y�7+chrr��Tj����ԓ|?���N����?��X0s�Q\��ɒ�	w,9cԃ�E���Jf�u=�bN�Ĭޔ�w��kx�"3/$��QUQ�1B�0�ڨ'��[m����%�B�ӄ��BS�x+�Ӊ̎��6��@wJ{Ncm�Hg�P뷇���!��OT@ɿ��,�X��HT�z��Ԃ�0�p� �C���1lu�Y��LC#V<j���%X��� �hT�1�n��qPA&4oBG�_��'<'�nu�j�n-8©F�6�R��:� w�V����P�v2L�B�Qj��Ϸ�4�F��ϙ���4�=;p�����9u����kR:J�!i�� ��y4�ď3� VR&W+��(7\)
⤢a^����
�=�Xa�@�"�m���q��հ:�Emb�ԋ!��R���0�.tq!�(�%�����ꋄ�th�@q^�$��MBK7C�P�/�+��?2a�
2@�.�uT2E�)��OZ�:�G"�h���O�.���,���	K��Q���I�Ȯ�߲A��NG�zo;��G#)E����� 	��j$b����"Ø;鬃�9�[�������s���!%^|"��>Z+�)�oA�����`0h�T�����+����l"S[����'�ev!OR��R��v��]ð�f���ԗ�!g�2�K܂�[�̟H[lK��k$���'霐�[Nz�.2qR'N��ĔBT|^�]Ng؁�0b��]�k��\��Y��(��@1�"�3�9�KA"���Y|>������F{�Ჟ+��ԃ�S,_>vJ�x���P{ �(6���H6��Ȥ{&�Q������;MX���g�|����[{�o�1�_�X��7�|���	r�׎)���G]R�GG���������X��"��@�K%=�MkIЬ"j
����}I�p$��=)}�v�|��7D��,�a����baL�����a���� E)����4�:+�I{����"n���g�Qk	�.�a�U7p�K�C�Ik�R6E�����D�d}��m���]����6h��io�)���AȖ�%�������:́h�[<��j�	[1�8���G�~�u��r@Ø����aCG�_���Upu�!�^7���&:>F@yT�8$�I���k?%@p�t���J��>���fh9[�E'� ��Uu8���p��I��Y��ɓ1��
�Ket�# �����1����Ҙ�S{��h����ѓ����θ��*B���+���D�{\�s��Һ�b^��E�Y* V�<cέR�<��dd,q9�I�ǘ���縮Q��������m����_��;������>x���_NsD�ḧhɧ��>��J�O<x�Fh��l����8���{�Et]W>�l�d�Q'��*�5ɤ��q'�0�w�ޱj��W�8�T��'a�R��;/���^�2�(��<�k�C���IP��C��q��a���85�����"[��������K;��Uv��=���Ϸ���_A��Y�耴�-��{03���8tȈl\�ڗ�;�zϞ�[2FWJ�e+u��訩�X��X��c��9cq�#Ѐt0(4�dI����:��a�u�i�C���2i=S>hH������믽�s�����G��T�u��*6�ߺh�/��gg4�j'�B�#� ʝ2�ʁ3���am�/���)SK��A�*�x�����������Vm��9�8�	��oWvq6֦5�/\�(RJ%�|����3h`tB��?�cٲe/�'��;w.B����ß������y��WJ?���Ej0�I_S��MCˆ����i��O<�L�/oQ�J��}���A%�Z��6������-����X���������yc����غm�i�T���%%W����c,_�ڱ�I�I#��+���?[�ֆQ^^�aƲ{R�K��۟�����ͩ�xm|e��\��ҷiVF�����]�x�0���RD�����0p������4���P<�h���'g��TTT������+��vdn�F�?��ڴƊ+��u���{6�yqq���Z�p�����k�0 �[RR�'��v��몪��2�O��hV��k+u]���a,)...�ƽ�o��*]-//�4�KZ�[%%%gfcs֭[W�u����cS4�Z�bŊe����p=�����ٸ���x�4�K[ƛ%%%����ُ���FO���n���0�b�0��������QB�eY"�YUU�@+��m�x�0�?�������o�ˆa��*�|cp�
\�	>?�F�=��ƮX��)]���c�_�|��0�m�16�������SQQ1����V�h4�+k�+W��K&���ceqq1-��s��kM�����8뮽�ھ�ؘ�k׎������0ލF�YɈܬ�]���0/..��{�O>י�yN+�������llNEE�����٭�h4zz6�v�Y]�/����=1p�@N_���˖-��,�W�b��|^66���bRee�V��v4=#k���뗴�Os0z(>��a����(�5��nݺ��n�z�g�e�UZZ���k�u]��3�@ �Ԁ?����(//�4��Z%�KJJ~��7f�ڵӪ���t�]����...�2���c�d���"]]�n��[�n��%kt]�x��?<=`��+~4�1�Y�Z峢�bzee�M�0�\��:g`nI����bN_��p�1�5M��CT���������0V��P�yXƲe˞�,����&�V����5�\��^Ɇn۴i��P(�m�T*�NYYY6�յ�a��y^E!��篺��~4�Ix¶��4z�r������|޲e˖�Y��DjL����Ҭ����� �G��~���k��u(>���X�d�R ��(�|��ʊalذa��͛gAZ:�&5�#G��e�ʲe�^�m�"�G\�OF���� V�\9'�J]o���ܹm�ϖ��e�Y�f͠>�����;��pgհa�f�0V�XQ��'I4k�����,���+'fk�o�sXy����Ζe��i�i���e��nݺm����ܹ�g�i�h��b�f�QG՘��w��A����$Ɇa4���U�=b�Z��6���Q%�H~��8�<�!ڃ�����92f,    IEND�B`�PK   7��X����(w  +�  /   images/42266fcd-641e-4cfa-a619-b442e1b7bf10.png�|wPSo�.,�X�( �KT����t�C(�;(�Ho��;�)���Mi���йI�}�9ws�Ν��a�	�d�k�{�g=�Zk�PMu�kT�Tה^>ע��(HAqf����贂��/�߽�s��0T �;s��39
��)��r@ϴթ��@�c��~^�Sy�m�?H�����@����&%`������;��Ɩ����*.#9οdC6��񕭖Ĉ�P��?Y³�T��^Ե�y���ݑb�ћ���������.{�?ާ��<��7o$�'������������g���+S�*�%+���9v�G���4t,�
�I�@A8=(��#�2ڑ���,�����u-��k�E�Cps%�%]-
ϐ��G]����[�?ffL��#"�yd����gP�==���U�c��\�}�?u�IN�OIIy����2�\̗�GOWW�����k;�-�YϤm4b����}��Y*��h�+�e��/�tP�i.Ӕ�����#�϶H�N"�ii�H=�).�%Z����\��� ӿ�F���N���/� t����Z��N_�~���ӝ�hY�4<<:w��Gxx8D�J����ML����#O��	A��ҥXm��k+���|�*�[c1s�Qf�C	���e����~s��oZ�/	�ǥ��{����������rw�b�0�C�t#>#�����p�1��|1�8��;����Y��h]�/��2����$�i̍=��3$�{����7�����ܩݖ�%��}W<2��ɔ��І������q-ԕ�k����[-����5(���Μ���h)� �7H榤 ._�m*�T9!)���l5Fl��gR���

�_#�tw�}�Y��>=:�9��)�_O����`m�q�vM��R��S�t�8���������*g2N=�-ʔ˲↩�ު7��ˊk�g���\�j��W�7,%����L��ض��h��	�m��V���O�����_�،����^�,�7�uKK���Ʌo�pq���Ù�� �5=4�����jɩDs�!�Yݜ�Y���b���nx�����s�g[o�3�6
����?��g���;wq[�X�|�.a�Kn����{�>p����z����� ԧk�Jo4c���;���P&÷W��\`⾻a�[�)��b����FFӃN����?���Ó@TA�����]��!��%����v��^�����K�j<��/e���nSI��{��T�o��x�{�:u��7��_vb��,":��5���,v��VKN�ê������xZ~��s^{�z9U5)de/�	bQ���UmB�Tc��H����Y���{�Ԯ����,7����;�c�����:a�i�R��I�2�^�2Jq���)++K�P�ـA�MIv9U�@����E��#�6]��8��GHڝ�X��t�1�A�ڏhy۱�7�!��8�|�jiG��:_)�t��o55i5��� �*����G����cXO��[�W�_���+?nph���k핻:i��p���5dɆz��W�@qX�����|�c묋]��S3���Ɇ�4�W�<�����kj�nrg�}�h����_t�N�D�=�[15�Ҭi���cm�^��v5*ύXe����U�u���)���)�lPCP������Cz�w;W��d�/:��+۾O{�����5Y@r�,l��פ��7jK(^0��'�^wm�k��r�������_^F�z�R����1�`@�{��^��ט�����ǻ� V4}��K�6�����cSͬp@:E׆Q�Z9N80~�P�NO�����V�� ��;~���#<	��e@ɮ� =���zo�W��L�SE�2"j_;��g,�m�+��i��grg>2�ޣ�dF��1��O]�l���&^�H ڨ�S/E=|He�/"�}�X�"kTލ#�R����l�:,c�
/��"M����٤Y:s�I6?����!P�#�9���ˢ�tE�Z���cu�ZV�L����'u�f�R��״�el�y�}x��?������"����c�MjMgϳ]sHL��=ҪaNO�
7& ??n��`@��F��F���r����W�{6�G"�8�snSѾH�f��1��4�a��#�'�0�u����/�.::�Z��R��6�
g��=!s|5���t{��2��R>���M�VZ����>�� �M<���=d!�b���ʐ}�����Q�4�_W~(-m�	�C/=�}U,����u�����=����Ҩ8'
oz83�y�z����H@�ˢ/��;�ALɩ|}��n��y�wꍑ�xj8�[���u�H�{��;��7���ԡq(��]v���X��ʺ�c��٦�B�^.ݸ��o��dO,��Ua٩�2���}br�3B ���&D�h���������G&�=^Z�@�C�[�o>&u�g�:V�9�m|���Ewt��Q��҅�b@�m-�6��l����}���&$�p��=�zq�<�:w��+ ��������[��'٥�+BZ%����h����i?
�>��ɷʮN
S�`Я� 1ܿ�� ����cޢ克�=AS�d�"qz��3�h���͹����̷M�,���_�<^%L{��"��l�A�/,v�,��_���M�8�"�f�2m�V6:���*�����3�))Qz�{�`��%�!�A�;D���G��c�w.�{�9���csz�7�.W��Y���;��B��`��zMp*�H�;F������t�?�s,�C���-e�z�A++-P�3����7XĪ���~�l�F��g\}���"���î��Q�l�Ԙ�T�kǇW�h^�����y%��13>bZ������C@oݼ5�$�cr��ks3{�Փ(��Z��dֹ�]Ѽ7�������Qe@���:�� ��/n+���	�����jXD]vxU�^�&�00>�ѹj?��۱�n����"7�l^ٙ�-�� "����+G�ϩ$|q������%-�e�� r��6#�U\�����m�F)G�e�*۵��*�u�Tc��#Ϻk�Ӵ��&^�E�g/��I��-F)1�z�����ί���c�|���vl@�]񍹢���1��a�e\����i�F`՛%�R.Փ��DȞUo���R�k�e����v��I�e�7��:��C�=D���{�f|yV��TM��.��E+���<m�P�)I\G���aoh�K�������L�U�n��/��Z�|U�&�[C��&�C�8��yǠ�t��H�
I���WSfn<�)�^�v�?�e�6�ļ��ã#���-|��D�1�I�3E�y�����D�NI+O.e;6U浺n�/ ck��S�XEt� �Ҽ��Xla�cf#@̾%N"Qע�MR7��^~�Qa����1���c�ny��TM��`lTZO����z��f���G�jȈm�,j��Y�)<e!ȵ��:���jDt{�e95K(���Q��z|��N�\T #�#�פ�q��s�޿ٸ�����Q(��߭�ފ�k_���=}�k�l���JҎ��M�U�D@��r��c��nk����2&���o˽o��K���<��4�ٳ��� /Х���߷e@�0�"�2���4�<@�G�� ��ؓ�0���Uȣ���v�EǨ.a��~�-]-D��`�fAL8�������aUr^s�B���R�a1?vv��3;6���x"�P�]�o{��풴�%78v�En�(]�8�y|�l�FP	�nfE�ǡ&ʵ}2N.�C���M�&���N$
z��
wq^0u=$�-�*l6	�n�lj<�o\��]�������c��&<j0��c,A�a��p�cٓR���#@M������up�7�f��@U��,J�|��I&L�W�S#3��ha�~��p�|��H1�2��݊��OivV4�`�D)g��8#��w�����}  �V� ���T�ݑr��F0}�������p�eW���=�: *�QK^�.ϖ��l6�G���(f�g
i���#�U���uNq��
ڱ{�Ƚ�ЃW^PG�D"T+�s���������2pD3��@��c͋l�]���b��T*�����߻��.�2#���"MRO^�4�o��hQҘ��";�x��͛j<C�,-m��0����m�+��9{���-֍����4%�Ia���J���Ƭ��,[���_f�lG��D�n%pYC|���>3Yg<9�Ey->CgO����|$�7����R��B:����ˋ���l���D��aV֗�Lf���?�����hd��@G��}o���������|k.��Z�����Dd�a����1< ���#���[:^�]5��h
ɨ�"V�����#��h�ɶ�AFTl_��«HQl�}�i;��o�m��j��b�N�z���Ѧ���t�2]�ĥ��r#x�J�H��*�V�.�EŉJo��߯,�����
�O���~�:h�ie���+�Q�1�Q�O��W��x��>Q��Y�����+�t����h�n��כB���k���M��(`1�n��P|�z�P��4=��H�}����)�	N����0#�8ݫބeob;YSܪ�q�JZ�}�o�⫔2�z���-����K�
wﰆ��	(�Vy)1�b����j?��E�h�V�q�����b�^,6�[XtVĈn���]��/O�#W~��:&�'��Q��J�(��qI����������1�µ|�e,��B�,g��lQ����6X�~�r�:!o۵��]��Q�o���@s@~��jC��V�l���̛�g6���v��LO�n�9F�y����c-���k �R��ŀ���b���ٴ��'��˶��3������������6f�2氿h�7Q5�ÊMbY���]�3�����Z��Q&�O��K�-��<�=!�BӁ m}ؚ]�l�r�\Ṛc:���
�D}N���U�>�<Z=���Ũ\��o�0�t 
@n�o���l����X����w�,����
�CӿPqs����$�Y�"�r��m4�G�r�����~=��ب~8�n��DU�x���/2j�<6�Y�	�GG��H�f�|�\��̇��ՠ���0Ҽ�.6�m!�����l�^m�$��}�Ww�9h���a��J��@�$���뼴��l�C�J����d/��e�>3?^) x���M��%52k.��t�\����t���kS���W ��F��2���DpR��T��'�d�p�f���� �e���a�g�O�յ�*�y���*i�w �^�(!k���x�TQ˚��$�}�8�]�L���L�+�GN!�RR`�����pۯ�5��qOn�Ϟ!F���b��>7��i���xShl0~В��D�Ȫ"���iR���;���15"�þ�(�u��*F+7�#H��:��CI����eF>ܺ�Q��e2T:XJ㿪Ljy.D�h��ujyW���kϛz��DX��Wo@�Lϝ)\x�{z,�U�B�VV�Ȗ!��`)�0C����9��ii( ++������uƙ��t�Qȃ�_��I;�Qna��\H��/���A�O{�9aX��9��(>�F>~|9U��`���Pv��7fs�'�2�7���.2TW�s>��D���d&�	�U�+d�o�{�(F�p��&9�1z��G#�cuĽ�%Es�OJ�E	o *٠F�۽�5a����r°M�h�}6A�P	`ץO�,�������(��m�Bxc]'m���W ���!���݃=�wD���U���Rm.�U"�5�_����WꇷP�g���[�<�Y��	�jg��i��Jtn�t�,��#%TO�h�
��h�˗��H-����`�_�L>�a6��rR!ő�6��|�����d������
R�tC骗#/H,떾Y	��Yב�Y��k_B��U����ի�)>>]�
T�X�@n�G
V<�t�!1��E��1:�?
��H�W��/W�z��%�/��&.&eyW�%(�!��)с#������f�
J�-) �8���Q�S�E.*2{`ݘz�"Ea�{x�bQy�h��J�os�q�(U�4��|�X���1��&c�U|���V��f�p����kJ'�ۻ��������>��܌�n{M4�B-|,��������Ђ���*�_}R�N��wG��C�b�E��A�?��m.�(�:/�X#
�c��I��B'���+����cb���&1�%=���n����kt����.Uf�uT&ڑ�c9�i�Y�]�7����������p�;,�C��:���* ��m�a4���� h?�s�.9 [�j	ix�v�k�Te�y൷���mU��S�L�8^�,�VS��Y��ky!sا~��}ڨCߢ��5@����#����f��hj�1��������O1l���蠓��L z��ge�����Ή�Is���~�bp߱��|A�Ll�՜nk�י[���:��z�㥶#����B���'�ʨ.m�`!%�M\����a��W�<��:��rH({A����Bv�1(k��vo�GI�I�,��U/�U ���#���ILl����&YE+{�|
'�ᰱ����2�Z�?�I���/�j	o"�f�[;n�|���Oײ:���4���kX�Tt'��B�BǵTs�` י�I��r�u�W��X֦�J�ݖ�T��$=�T�,{���a�WT���5�'O��J�������\M_iY�9�}|���G�9=��M�\���hw�p��������զ�	B��4_�5��� ���N#r��'UoS�RP�b����!��cs/���m���T���G���zz����[�}�&g�v��c�P��Gc�e�C�y� 7e�t�<���!� ?~��5�q�>�zF���{P������h5ns�0��h�I@��ߝ��p�g  e�7��~[�U�,������F��#���j��0����ְp�2ouD:1p�o+�i�3zܰ�Bc�G�h��e+*�f$!_��Gv@��ъ����"�Y�:�O��﨨��|����3#�c���Q��{�Zll,�fny�	|Ks�	����+��&1�e�j���J=V����;�,F_�FLnBQ�"�{o_wԻ�y!���-)S��s1�|��39IMy`�n��G�$]IyT_w��Y���Ⱥ��H�hi%�7\�5�������i�u1��-+�,��Mx�1��`y<��*q�M����3#w���6�Bk�zm��A3��V�ۚ��-��Nn��W��|/�)9�Z�����C-�] :E�b0���S�Htq�G�ʽ�Ws��yTB=��J�Z�� �<D|�o�Wqp�Q�wo�Ņw�Fvk��BO$� �珎y��ER>��z��^n��=`6�W�\gU�ufZV��˅��g}�ɖ����W�����c�����isv����fdqQ� U�J��V�����t����ƫ
4Gp��Hy7�G��!��zX���0�Y�e��ڬ�	�̭&]�h�^wo��ʳAAy>�Y\�D��ڧ��=�?�6d�5�?s�E��&c!��F�u����ʝfա����{S�W�i�c�K��]�������j���kG�5�B�S�\}B�~���(�Ư:�[����%%��������6�5W��.]���5���먥��׮�W�����]�P�R�j��t�]��V�|Y8Zjx�~�F�x��A�?��F.�}s�o�5���<��⡫��K{���Q����f2�dO��f�O��)�M���X�Vs$7��|���QN% �)��d�@;����i�1c��2tD�6G��ԏ��s�z�j�ݺ�Ҿ\�y���(��Ħ�"�:Q�Q���3�^1��gy�^�vu8����E���?�%�Q ��D�29(�*��o���f��yJɣ�B���o�~���RT��0H_8���=n#F�NN0%��
D�x�ey�~���e%�V�T��;����tk�2����-��i��IhǣT5�7ۘ ���8Ul�4��؍-�é#8��Z㚄x���<.��C�S,�	�Y�[�r���X�W��I�9^�7 2�v�=�j�oθ\��w �s���򄋠z���$���`S���hIZ��}&�����'�i:�	_;�p�p�o��~�wQW R��}�[{���?��1��2B��Oq�&���PIk���ٛ� h+�9Yp��]m��{byΑJ��O1�c��ʼ�� ��w�VF��Ei�&��{�#���4�Qq�"uO�x*􅍾NG.�\��<��IR������*}_U��  �f���=/�N|�lF<3���O�Z,����s|���q���`nC��`EoU���C���I����P5X�/��K��6h��nhn�_�f����H}�ciO�����aCe���aM	E�Hk���l-	����"�ᾡ�-t�O�fc��Bc?�Y1�s���9����V����)T^b� �UVd�pS�o���ߘ��%����ZT�����qF>����6������-הS$�NIrق4�q�5��D^�6��B�R+��/��G���	�}u���r���X�P���V�C�� K��È�x'5.�KN]�F��_o���C�ɪ�<��SgڃT�X�&bY�n� /?�>�97�d>�ڶ9s�䌗/O3��&74�K�J��'�q uf�6�CO�I&NF��o�3d_/��E"��wxde��t'^�T�nD��&�^����|}���åo��W��_��1���Mf�z�y���ըX���$7E��������%^�i����I2C�>��04�2V���wa;� A$'#pA�1�%�n�%cz���...�t��<����x\���1�5/8vr���E�92>�t���.��y�~�{�,��)LO`�����JLT�ZKH�㱾�<v���!�J܀a��(x3w%��kz �ziZ��Z�u��s�B�JC��z��_bq]�3��=�5!$�(�;��#tx�z�n�q�D5�ʝ�J�#����>�/l��������$-kT�L�@Ña���)LhAQ��=x������|S�x�ɖ�%��)?~���{��A����T-�m�Y#y���$ӗk���ǍwD�8�Ŧ�	�	�j����<<�+�RV�&�ȒZ|�}z�fů��N��fa#��i�o�o��xab��z<ӌӹ|���W.z��l���Uq���к�!M0����	tyC�v���ZL�yo']�]?����2.�|�R��&7�V�����"�q=;�K������zy[˂��o����|�G��yǇ@r�1	���1�)�5��9
�� J��?��T���v�9�$�mNw����l�+Ýֻ��p"�)����0>��Q����a��qL��/��g(���y*H�(6��0d�>5
B��?�
u}%���i�a{���{0O��X�t$�R�P�|��;�m����ڕILO���Ui?}��H�tR��\�B�,Vc�+m0 �f�}���~�"c�&�M��a�\��8��t���\��.v�ޖ�Tvq'�ơ
n��8zv�w� t@;6�cO�p:v�l.�A�̼ݫ�|2�VL|�[Q��ή�<"�@�����P=�s�V�"�)����b֭���s-��:i	�2��.e�|��E��"W��̂i֯�׾��hy&��/�	h�2�U�>�X���d�z����a����XR���֘�,���;^���\��m!�WF���ޘ	�
���%q%�0r��tGm�
�V
�en8ޞ������o�J49�M���=�����-rl��k�U���<�	w:V8O�/�:ױKtq){��B.��_h	�s��܌�;^>�H�XM�	�o��IHS�)�4�M�'ϋ�U�{۳���ȃ	���'��, �=Ó���_�ZѺ�r�@R*:�"��K����Z����pX�ŏ�Z����؋�D��ߦ��2�ΔM�AьdC��m�]�vVl`�YMNw�I��z��P����dE0�}\��[��~>�Yz���$�ůӞ��{"<�ə)Ӆ�K��#~����^"DF�����7�+h��2�뭻�,k��wƟ��
����5�ϔ*�*���s�"�Z���X��l�ӑ�so�"PCv#�3�D����s�d�Ulr]���㿤)�7��N6�%YYOߜSIYvcv*V~(i�}��h��6~L9�M>q��9��b��G��4�>����3�)7��m���a�e��=^S�G������ix�qL=h�L�wN�8 y���i���e�
<�K-��K�lpn� ƯQHR���ML��8E|b�*a7�{݇�Gc)Q�	�ņ����$Q�9�09\ ٵZ\x}Cj�z�.6����ؤ>S��:|1f�����k���3*&��I��	�8}���7��ٰxSs�2�2���C�L��H�wwףb���0+#�Z�ۧ9a��+Z����o"��5�5*�"b������f=�B���~�F|{����UaF��[�)Ά����6�Ձ^��?�Y�?�oܖ��W�2��M~F��ZZ��a�e��ɝ%U�Id�x���~�"z�A��<�I�S��3mi?QFcNZ��E;2P��Y���j��JC�����f�)V!�O�Y����Xy�������N�i���$/}ל���l����7�댩���][�1!�y����Sߪ �03nlҜ1�6���09�V�L
xX��o�=�{\�����ڈd���s=r2d ;��q�Q$�y\n,�GS1�����S�F}�(�l�qT�ʗ����Q ��2�Z+��y�`MH	n�"ۙ�`K�O/�����8o���\�����S�V�/��{�U����.r�T�	9&�5�D�¯�݊'��[�D��
���j��>�IHX!���lS����5��L�8X��c�B�F���6���
��9wJ��=$ZDFX� 2�:����!�sW�m�9�o3>"���o�=���	�	Rm�5�Bu���"V!�G�ˬڡQa�T�B.���l�Ge�aɬC�P0��XF�o�ҩ�۫��q��L�۠�r�-��wQv�;�2���s(U���)��� A�y5�����p3�5Lڛ��\�~�c-mTB$�Z_@���p���p�����}�-������|F�jG���%�"�%���>��췦
�Z�g�=P^�LFu6j�Q��r���)��/� �3��U��G��XR_(���B.��ٕ��$2����<U��V��j��	ҭР�N�kl��}��5JF����ųU���0U&	�u��TǀQW��Ӥ8�=�d��Fנ�����ki	�mM��*AZ{�)�������e�r�LC��������Nny���	=����ņ��4_���Z]���dZ�����따ߖ+׋Y����PQU����<H-�+Ź�ǰ��ɻ�o�Z���ex[����������֪2��5 �/��SV�����{Ǒ*���)��pSJ"�xZ�٦<��6}�}�w�^
u�c�O���a��:>]fn�����A.ۨĦ�Q���ve"�םS���J�T����N2��dʹo�r ����5�b�I��	cT�!5�����3%UV����s�i\�\��:$�4�=iP1L����ã3,cEĲ1#"�ɳ����j�쥢�q�Q�}	�v,0���X�F��+������â�����@O�f���k�Q�2M�h&7]_� �O�k!Lq^���ĥzM�t� �����O�~0�Iʹ�ג\!����;>3C�A�Р�$r>�_'���U=���4����*��AU'o\�\)�`>�v8�U'�C{�=I�M˶�k�i��?��x!�O��F��,���Ϗ���L�&�����➢�9jUj��D!n�{�#��)?�;���rΗ��}���[q�*_n4��E�ˡ����{�����OTo ]�Tw<EK������!��I�Ï���U��w�E&`����U��/@�Nï.��n����5��!�&H����t{㑼�osX~k�c���9r�#���TF=L�A���O]�5����*�/Q��7ʈYŇܯp��0�B�����_�s�^k�J�+��%��w�tEʄG��=���+;�r�	l���F`������ve�Ʈ����{���梚=�-�r)�RLO6��2�?w�Cdh��e�-M���[�N�  �͵�P7��5*j����P�����<|w��."�T�?!�
��[�KBnB>��N3�"�D���(��_�S��~��y��8<�Պ�?���!�h"X1z�; ���f�\�TuEX=Ó5pzuGw!�N�$��]ɤZ����0��'km�!��Bm���O ���L��� 鎺���.��x-�u��%4忹(
C�.L�P��5�hJʓ��� ���a�F�Dݦ����!���,��:��_��v1��+���,_H��%��-�{#/�����I1:=���[�N������T����jkx�}�a����" k�r�u���/��/�"�G\���L7.���\O���
{���R3�jE6쳶}���S�c_�c�6��L$Iח�C�ܮU/�j&�x]qk�SH#6Rp��`��x&<�,���AN�I&���MM��V#Ҁ��v姱^����ɲ��
e�_�h�A�,`���b1���A��k��,���4��{�5� �	+ߞ��v�=ĜkhepY�>���^�ا�G0�P���/ז&���?�qŜL�0T�B�7�iv�9��k�����6��߾rח�:*\�,�,��
jh�xݦ�����9 ���d��Ŀ�H����Y�耓x2�&�ʅa�mKn�L��ϗrA�Qb�}5����ߦJ�r������8�W���U�w�ϯO�4��$��=���{�u�
hF.�ɜ��_�U�L�Z,2��g0�Oא�ڈ��tE�p��ڈ�����*|Ο�jS�םS(�����A;$[<��_ s���i��^���05*wl>�u��Ĕ�<����n�,����@�lb6n/E���ma'�m ���`�u�飽D�����kk�I�:����V1K�(�c�
�RH="�d���1��M�����Ot���]�⣵��Q}��I�=���-�lפZ_�0)��Sc����8���Iv6gG�G\v[�3���� �Tq>���x���c��Eg����7�U�dPҼ�'2>e�I��Ti�=��j��?O�"�H�OK��p(t����iD��D���΂N8�C����/{α�Po;
Yv�[eķ�a��������Bk�� !��0h �����sx��m�0�0c�y�c�fO���|�0�]�)>ZJtW?1�؟-O��wux<ҟ#���&E��P~��.?��2�Y.�U(yc�\.�����R<5�Σ������Q���s��xD_�0�T���Ym`�OE������fuy���}L��WF!���vN�q^��U�ׁ��%�$s��>xj��18��2� &��h�u�	����ohk���:l7ЯE(��̒�l�L�c��n����	T����'�������dS0s�Q�B@nr��s
�Ew��05�,�v���Gt2os스FИ�� K\���`kC��b�eP)+S��"�Hҝ'ͫS�Ȏ�<�%�h�y�Qn�ާ2��C�:�A�q�R�~��L�ƭ�4�<2���l׳�'���_A��2��XL�ɲ/�h�?U4uze�f�˶��6��v�q�y�<�r��q��ј@Bu2����_+���3ʤ���g䌳���t�Wj�|���&N83S����އ��DJ�W�sJG��\,��U���o�")�@2�~yU�K���ޑ�g $>��q�q8M/��d#q�u^c2�kS�3xX���"0h�(���343�(��J��
Wmܢ^zc��|�]�b�)Կ�+��%D�f��D�;�(����jY*��gm�,�[�U���m7�6|5��<]�5�]�ȷ}�������~�െ]JX���ր.:��f5o�F\�f�&�m,U^����f�gGނ�n<N��"5��R��D�W��19���U�#f�h�,.^!l	�p�Y*��Q~���S��X��4g�\���&x~7��o�ᵨ5��QcHuO���w_O@/���Y��� 9~szL�"ߞ#��L�~}��#c~L�X�/eז%2b�&w�&yM��7^��̘s��/{[:gE�io�O�#k$Zb��:Z<��}��	-�r�U�z�ח�|w�����p0�V^�IL=�rJ����?��ͱ��]g�I���&��%$���D���@��Z��fK�|�)	��a��`�O�0�`�t\�CGs�q$�����x����-=�m�}-}qY�~�^G�=Z�Z�]q�<.J	�j$"��\-?H� 2L`���p�����'ہ�=w���
@%�*�G��0���y�³�$ΰq�ּm���wB�����כ��醩M�_ۙ�=QG��� 0�lP�@�%�m>s�u���'��<� M(�?{n~6ߵ.�]��0_���aT�҇�_-R�ɾ�Fλ��l?�¨Fd^�;�uTZ'=��,����E�S����1<�o�D�������F7X�N�	k%kuz�!�^W�=�P�S��ϗO��(�2��� {}Y3:s�M����8��q��*��/��y�>�f����y�)��2��|yvq�)kJ?>��
���˹�ʿ-N=��餋|n7ļkH��u(�V(�{�α�.2�a�ٳ��Tf)ǽc ���ǖ�G�RdD��n}���^��{R鱧/@9�5�-x��[ A�4���(hC�Cb��D�<1�Gmɐ���)�T�����5*!�rci�������m���**�9�E����b���0B��n關��z7�Q��*KY��i'�s�]��!
#S�v��#������8�.��B�8]�h�MR����*���0���.r�ܔCAqz�Z���z��g�,[wY|g�(�U_��* dܸ���>���mcy.%V��+����?s���)�Ғ����0}��G��yO���E��\3V��zҦVZ7��f���V��}2����
��������u��.�
���HX�
��F<�t��|���BIm$6�t�"�?��Ms�:������W�G�3r��14��(g�kH�+��Wk^�*l��?�{��3��X���n�ct�y�ON>�O��EO��R�;Ғna!Mǐɍs���c1
��{JI�G���k�K�I���"�����~?Q�5���J�����e��'.ߤ��i�O��� �?92� ]����}���_�Sx]��0�#Ht����П��`���϶�^�5��[xL<i�yj)cu�p�L���݈j0]���j;$�����w�?(��|�]aSl�ȣ�Ba7���ԧ'���3��`'���V�j�Y��c�*y"��qw3��+�������ޮBA��ŅBt_i9hF3g�תʄ�	%_I�?�����<,���[ە�0ბ %�E^l&�}�ph�J���2�YG������^�<ˣeL&R�_k�o���c9��vC���f��x���LBZ;���D<7�J�ߏT[�6�Gm���8T��T�����R(�h��G�7><,����䄻�ў�mg?�@%n�4�zL�Ov���D.v%�~�4og�w��6�.2G�p�B��uS����1�T;��������ӜY�ڸ��5�X��Q
��^�d�)���x7n�K����(�Бi̬�/����L�m��yBɍt� ��&�� �;���d�%�VӚDq���O�Ϣ�}�ISk��K�JH>�]B��U-��!��٭�&>�1O�Q���.�����CC	��C�	X��D�f�EG��� B��87z�V��W�D��x��9p�a��rӇ�2�9N����6�����Oψ����|`r?�x���+C
T�S3}d�{�����3�8ZZ&?s�q��"��u���{���g9OTym񘛸����2�I@65,��^��[R�]n���Z�'��;��u���b��qد�����8� �
�aL��L��g��̱�o����{�����[�<U�"�B���/l����	}��_Iy\�?�{�;_�����--A�Z�u����yb�m��0M\ ��p�^���	�4�vDv�{Sڲ�n�xLs�8`�qS�UR����T��Q��̟�U,h�7�Θ�̹[O?�Z�Z��3(�"fwoDm�����xǡ�m�h����X�a�8OS�	?�����K'���;�|t{�gp�e���c�uXW���)��l�z��p����I�}\�1�=k�uʤ�04���m��%�
�*u��1q+UE�s�'p�^Wn=�������`/��fEl���xuE_��,E��w�`�4n�2_�4g�>���P�ڥDg��i��R]�*nT����o"+�u�f����H��@��ل�Z���F��v5�v�H���1sB�Q�1��V}s��Қ�׵㭹z5^����\�#k��e���ȩ@��}8�f�I�"fF���������+�[�n_�;},�`�����KEj�O 4z�*<���X�A���झ�ݝ{��ÂO ��F�KaOY>3���>��5����QBb���AQj^����ޣn����l�z����L`N;��U�KĢ�k�
���Ku��RT�g�)͏�!��i޾�sT�O'��#��G#����i
O��7�@5�N[�)�v���=���On5{n&N��R�}Pי��=&A�7�ϭ���#�H�|�f�N�I&@�T�����
7��D���fĴ�_)G���w���������jrk����9r�RP�IWQ�HD�(�!���L�  ]�=jh�A�H-!t1�B�y8缳������o֚�<���.�u������PQ�
7g��D�������B�_g��j[��qB���!�5y�/�g�U�P�˃��[4�����Y����ṯ��F�X3D�����n��e*V��l���!�<<'C}�fg%� ����� p� �P��^�B)j�?��\��\������|����n�{чK�Ȑ����x�Jն*$������rG��̢z�8�Qmk�{�9vj�sY��k�Վ}����o��U�Ϲ`1/��<�Fv�W�cY���ܹ�������>~���e<W�~�`�^=�U=�W�D�M�;3���*� �x��K_��C�4������uӧ(�6o�zf29�6֎膿�� �9��M�z`�!#�9�������}B՚��,C���Q���c��)|c���}ҫ�g��U�Q�9^C]/R�U�������s�ŎUx��r���pG�A�������w��ß�~g��vLTF�y���5²!��-6�b���1���x�&p\�I�{�^�_x�?��t돤�҅H��H��~�wl�|vU>�9�k���xB����e�'4<���7vҵ|3ɸs_���w|��W�#�UM�l��Jl��Q�	��wi��x�u?�L<Z���6�'���"�Lx�D��Q�`KˇO�!,�X�>h}_��LC�j�ّ�֑Y�$(��!���t�"*��_��SPyֹ3���f�.���;əp@LWfݪ��0p7�u��撥�Wf�Y�aN��X�]܀V�F�4,9�?�
�.�d{����&����i���Q�M�U܄M ���Ym>�W?����9�Ӵ�k]��u�7�J�0��"'~$X��t��K�V}�JR���]b�2�3��Jd:g���r���k�d]��Ĕ�ڎ�wͽ�k��n@��b_���w �W��×1 p������M�������GL� ����t@-���{j|!���e�\�8�48�����Քj�<�/,Y�K��r�̖tz$�H4���L�����M�+`"�����S;�4����ؤ���4٩8�k�&����ڈ`����@6���3����s��[WDl�ȝ3l���t�8�o&��Lt��Pa羥Z˕A�H��N:u���\ bS����v�͎�>����ۏr�U2��R%o���d�b��czS�U�ě1�L����b�r*u���c� ��%�q�!
�٬AGB4YU�t�4�RZMw�j	ݻ�"G?��2|�����Z��XblǺܝ|���I�-�9������8��ae���m�^D�=�q�a9{�/'x$6t��5��Лte5\���o�!g�[ف����Gt�ֵ¯0�g�h�o���ܙ1�;[���{!9a��y7��+E�/�eG��, [U�V6y&�J�Mc�eOՐ}̋��Y!2GBE��^&�]u�m�a�7 �/��]�5��8���m�4�� ���������e￤���a���c)�Y	
�O��du��S �΍KI�uA)�y�P���^��S�VqZ���l[�&�:�j��T�,�$���5IH���9p���g��me�r�]aW�y���Qq�͝R�U/��T��|_���q��\?�'y�VZTl�,)*q���.�����yK0F�����`4�I�@~�s<�
���2Z���Um���0!ſ8����!Yo_��"��`OQ��D��g��h��.�4R.1~�t�ė1V��nݕP}�9z��)xI'�"GĨ��"h5��Ǩ@�[�z��$�d5`�Ĝ~��ͫX����ʇ١�������S�A��6��&��}�}z��A8ܣ�D1˛����q� �M�S�ZFV��ؾ��%�b%��6:+7��`�o��Z �	�.�y�U!~��D�ݵz_�������7�8�Q�����]m�ryq�e���gu+�	 (d\�F��u������K�����ɵD�m�S�6y$���I�Y����P�6`��}ӷ�k=�c����]�/|���Td*�"8�}�I���*/��,[�"l�槅3����o�",c��#m(��l0��(ON��C5���ww-�}�{�ez{(��wX.1���	\��LXU""�#�oʇ��x���b����W> �/wa+r�K�4b�ןD�m��:J���MP�m������7�Gه��N��T��#e=C���Z)��&_4jX/�Y��3�l�z��r����V��E?�~&���y-R
������)�q�
�0*`j~��/�q��LZ����&4Mp&��gi�n��!M���/�"�l�[̺2�ݷc�)?��P+�q����h�S������j&�o��{l��ec:,��ߔX�����AK�6���rG[�?Lq^P@��m�Ȅ��ލlEo�fb޸�)hi��ƪ�7�ݚ��gn�Z) yHk�_������X�E��_���s{ a_%�T`׳W5?Z}.�C;xD�x����^��ʀ���8�!�CV=~j��EJ�]Aw;����~�]�F�����>�vq�1� HEHY%V5�z�P혡�Y�|�^}?PӍ5ISpU���ѵ�6E_j]��͚���-
�Pu�u=1�3�m@Ц�WWn-Mx|��"�7_��y��ј�DU6���N�Ho�m�����q�>�Y�c�6�ޒ�t���w��4�1�K��f��zӸ���@˴�۩2�?��@im�Sj����Yr��c�D��T�by8�(��?��q�:�!�˾��42��TSҔ8�cI{�P0k����_� �M�H�
�g7l%Q��jw��:Y[�.<%�j��"kSd,%�6D\F��S��h���e5�}k	���3�i����S��HA����fϰ9àt�y㣭��"�89���:kn_;)k�s�<�紷O�(nbV!�̖�*�E�"� *����i�6O���o��D��4H<�.N�޹��ؠ.��e�N˵�F1J�1O.�_�U& 2)Fc��(�бґ�1 ��3��fF���$���d�������gJl �t�h�/ݴ�O�,sPvz�'/{�������U�ݠ�H��A8��P���8���)K�{��i8i��Ȃ��6s�AZ�u�#X�7����J-Q�Ɨ{U~���v'!z�n ����I���*B�i� y _�&)�G��/U��cs}�S�∴o4�5	,�R�\!}Z ��^��u�����h�I��X������h��4��H���gW�on'9�GHH�+gv�"S��J�{��l?�YM]�]	��&ܱ����������#�:�r���:�e��R�P*�zU���5��OV�g���jZ] ��F[�rFv�7�,���-��KM����%��5 �
���K~_��ji��F��F�q�jW~�c��G#r�q�g��%�e��A������`�i�
�s�]�`X�t~������ss� �q')�*�j�~z�,%%S%��^5���.5�+�`}+����V�~�G��vXJ����L�$2<)��k�>�t�2�����ͥ\i�#4|z�^<R�8*�n��l��]�U�1,�l���Q�̠{Òr�Gkבw���u�
a��b����R4��̪�.��8�*�h�7���L����q@���G>��ןt�a�W���9�'�oC�E{F	Hx2��:���_���RH�rW�j����Z���O>V�\
�q��_�=�.x��*{=?��0����[W��5�9���H:N�BR�1�ɪ�j�cb�+�y A��t�9���U
 0Y?Z��h���m� o_���� қkv�����GK��1�ha�3Ո�jK�������u]�e��s���y�t��Lx��(���ˏ�,D�rܪ,O'?>�si �3UE5�&���~G8��a5��4�ޠG�Gq�:���˶V՜��Դ�G�����'S����X�����2`T��^6��~���=qK;}���Yg�u���3T-UM+��9h��|e����n���A���|-��m�;�Í�����9��l�M�����x��ԟF�h�r�M��/�p!�19?�^)*��b?�(.
8{����U���<5|+��x���덵�I�VX��@����dSz�����ኀx���A�j1�z. (`�>X~_E>e5cI$֋b]�b9MՑD��n9l>��� �t��AQ���r�W��	��o��.%�k���]�m��ț��Q$��������<����w�e]|K�Ҋ&e�՟�^}}���5�,F�rUHVm6>g�8�ԑ �t_�U�[�H��5|��6F�5�I�p@�y�/�ʗ0��G����8G��n6/U�FW���S�&(	��1 �YTX��L�ϝ7� ����1n�Yt�A����#f�p.q���;!��AiOȀ��ٷ>�,�5�s�5WxT�Z+?�=�B2�R��:�؝)u��o�}�)�;��z�-�/caN�]��� ��(a��]�Q7��5�%�2�8|��Qz���<�SvV%�:Xp/wk^�4�XwE[��!5�O�>}23��,�.�;����/��!���\o��hm`�Q��)����uN�u,�d�GެdH���|T񷃇7�`A.�������4)@�}�ʣ���G	�K	a�ϼ��r�9�8-*
����{Du9~2�{����L8��}�H
>?��t�ݣ?���������C�$1;��t�cS��@��puiO��B,�f���D��YP�-�aIY��xJ�5)^.S6�Z�8�S��;��^;��t"�<�M]��"Fȗ@��A+mΨ�_��9��5z+}�����˾�c/��:�w��D�e��r��-�䉷���{8@�}�ٓ�fT�LͭbZA9���	s-�Vl@���I3:Py�����w���Uu�HGX:��ݤD�T���j�@��k�Ҧ�ܠ����Z���C�9�vD�Ļ�S�=8W|����<��J�p������gN������~���M�^4
Z��j�4J4Xo�����f�7F��߭�;�8������	p��&ݪ�Uό��Z ?-��[�i2�=0�d����#:@:L`������&iӤ�O"�nk�$��+�gm;����0(\�I	[{;����2L�9�b0b��<3wm�Xm��	���8��� `��1���8���z���F��i�MjYH5�G��j=��J�7",����-,�ļ�ӌji�%�,!n��XTc����F��ru� zg�*Lb�#Ζ:+��!g�W3%bVu{�T/�d�/:�S���Y�E@��
�.4�����mJ�iI�Y� f��
^��+�6ؖх֛�b��]Z���$�(��n���(���ͫ^nZ���\�G���=��ńU|�l�{�`յ�}�"��̞�gV�8�{�k/�8��6�02���y-�$�'�a�V|.#5��֥�[u�q�%�FP��d�^�y��q�;�Q�0��?&��D_
8��'~��Z#qc!f`|U��&rasƀ��BC��K�'�ۚ��f��N�Y���4�Go��7��Ü�k�o����p@w	���6��ix�nwF�i�ـ�Z ��Htf�>�I����ގʻb%�����
��9�%�#����ez��I�u򨆋]��}  iK��6q�y�4R�Y[���հ�<�����1l`���8�-��!v���I�����CG�v�҈\]���|-��f��am����o�B��
��]��,˻w�W��՚���M�r7(4����-	Q�_>ӡֹ����GNq��;�T�����w�����T�;1�!��Fak���4��L4��U��m�H:���.b?���-��fK�3<{sĮ)�>p���^��'.j��xwb���
��k�á\�i��[�
�|
u��qaW�H�B��q�t�m��Etx�pdk��ڼ�X�h^�u��	��#�x����QK|��J]t}Q�l��a���=�^w�_����J����C*;� ��[�3>d�k���p:�c�W�E�Q��ǋ^z9&���T�nHF�u$�(�)xk����ҫ��������UO��pY�.�����o0��%C��{+�p��n�TV���7��l�Í!?1�$�׎�ey>T�S&�7Y�>�%o_&_d�K=�z��S��Q�y>$f���kw�9��}41�A"G#�1����:�4J��z��烏��������gyM��� ���8'�l�r���e��<�N�>?FI��2��
��/|3<3����TZ���p�Ƞ��B�2"�Mػ�X�3�љ��Y�h�?'ez�kpa��� �bgA+Ymj=�6��^=�O ����.�k�??z��F�-���0SY[�jg�}��ѥ�gU�����&�P�+�~�Z�Dv@��=���K}Pc�B�����Ŗ��{mˤ���O�7h�	���f7�3 |���V�(�O��%���˛N���=�����~!�B>�)�,����4�!-d-�rc3�Aߥ���)��r���_Ы��Xg�}p�˷W�EFE!�_�����<`��^#PVu8�<��T������i��3�4�9���Zqŋ���L�9�vHi�!Þ���Ĳ	�<^jC�4
�9S���Ɇ`�����7���@�߿�����j׌�CCr��w��B�q���+�}�Ϻ2��<	,��)[�⡲Gk����k��s�XD��J��X�\���P��"�w��k��pD�/�uE����?TR�ȇ�߷�{~��p�	8`N��� �o�b�ƍ����u���]�jG�z��v@P�][�~���`�B����%v�`��+�x����t^5�k{c�ng�e��k�$��4V[���K��I.o�<�	���(J���.�/�IA�b�΍��e��,޲��t��Q["��\��?�b�'�{��4JD:���&}�vr/�V$��l�i��4/����OZ���}q�k�l��[2�	-�%$�1�w�6`���uo��
��g�q�- ��ȁu�KM�үF�k7���3Gk���O�MT�h�p+��?���?Q�D-ts9�5�'v$�s�;�dἥ��>uc��߄�G�H����O��q��Y��.v$z17�'���E�/Yug!���
f�`i?���bop��[��9"Uoc�GWp���}��ڢ6,�Pw���ٵ3�(�.~#���݈/�o��V�����2l=ve��I���x�4+���9�M�?}�ґMoZj��|�Y���+�� -�Z��n@ ?���q�^oC�b9VUzf��\������������B =t����b�S~Z�yqFƓy�������ϑu���O�:�O�Q&Q�<~}�?4ĩwڄ�zo�/_��O��|ރGm���͑�ʏ�C,�����ٛ��܉�^��ޠ��g/]zP� � �㠂���_�;Q퉒R�ݮ���R�	{��Kμ9�q[�Yx[�/�W�����Aq���+�o��4��;5}��222	�����յIxg������6K��GQ��q�3M=ٓkfY��^m��\�x��F�\���䵽y%��J����,Ǳ�����,Q6ɵ>��E��<���E1���|&�p"���|22WE�8�8�ۤ޲^y�x��K�|�m�t��Ƃ:3CR�<����������"���JC�P��pxc��aj�<{d�*���#��0*�s(8��u��y:M� I���mK��=o*�Z ���0��v����&1�m��6
��K�4�������
D�y�T2���n6?��Og���;h���\�����%�0�leصk�g�|ʎC q38,W�<�y��]�~���:'{�pE& J�� wB$=��(�������)vw�g�̌U ��^�2�+q8q� j��G�o��c���W]ʱ��gv!M��;��W�(�x��Z�L94����y�Ov�E9���'�׋���w݇��J�����B����A�-X� ��iɑJ�֝X���c�nk1;�-]����㋡	n��B���E_/�!��Ԟn�Ihf�M.	 � �>(�ݕHP<Lq��͐���7|c�s���"�����U�o]�^���$� ���3=n5�L�`��#��+�oTX���E�%)��P4NV�%{[.�o�=��'�6�oE��R#vC��C"�\���0JS�8�K���
�O��f�y`Hy�����^��&n�g�_癮��IՋ��y�(.z��\6*���Lz	��=��m�2<@&�9? ���51�i�ݔ�k�6�1��Z '�脮�M���.�<��i���47�a[���5�<�C�9حI�ەh�3�� �� +9C ��۫=Q�0{?���&��3I�V��[��#8��g�@6��*6�Z�'2Zqۋ��	11`�}��i/?m�^���Gv�̍���{����0f�U��-���f*:�(�Hr,ȇ��ùb�,��L�P9p��Rpu�/"���L\�έ۷ۜ;'_�@o�@��{��fl$/"E�t��~�^7��*`#�J
_���Ͼ��P�G�e�l.D/�~I��މ���<Wp��M���I��eO2,�ee":��ζ�v"$w��J8c��!K��Ke�!��?	�g���E�Ԭ�@�>��w�R�su��)�פ��\��&%K���~�[��+KA���l o:���k^ `�,:�(�JP��`��{�X�t�w�9�7G:��(AZ��l���[kY>Һ�Uqq�1%D�����_�����i���
�.C���׼���Y�&W��B�:|� A�X�4m�:us:=pqC�8+G�^��t�y�s�7F5������m@9o���۹g�z~�kgkx�Yu�ʽ�ۍ7Ϭ�I){�Q\5��r�ح�}���4SM�^���;�e����E���fi���f8�z?�	��=Z�D<z���YJ�s�����໒,@��7/��UD���+ N�{V�]��r����/}Ț�Id#��?o�ޓ�s]��O�u��V��:���@�*��S��	�,=��f�G"����p�p���˃�X���"����=EM��~�/C��~8J�����Fk�u3�#��x�3Tl�DP�w���"ӅW��s��pĭ�ij�^5��%b?�/��1v��C	)0�ƒ3|[ůP���#�&��.aC;���;��s�k�3��m[#PƐ�Ə��UٯV�>�ǘ?�d���/̣�2�u���1��[^'�>����`|��^��-���v5Z�k>�3��>�����'&�2�b5g���3��c�)m�Dq� ��W�ϫ�kl|���6��-С^֍��[w
kIA��|�`1R't�#8z���H>�#��o�Z3vL�����7�BXz5�1���ꍲ|��hH��o��i
P/��wN��������3cf�����T�o���
�?۬�5?�t�)V�1*d->��
�g����z?:�59!��N�>�{�k�۟o�`�O*�|:�
@>���K���_�������/RJ(���h����@.����ɡ��6V���G[���(P�����t ���^����h�|�������e�/�5��Ĝ��*{]����/�돏,p��c�N����BZ�S�k����'vDT�Xy~�I*��v�晀@;�H�MR�t}U��'&"-L#�����(!} ,vy�q���Q� �q��h��g�X�N�ȉ�j�C_��n����Z���*e�G����g_���O�\Їz��>P
�R�Kw���|D��ˣ�j&@L���V��;�4� �� �+^|�J��+��$9KGwA�F[�����H�y��m]�1M:v�p4��zg���̗6���@�㒳{ ��*^�H�,;hr����7톮�?9��!`�nI��<��sl0B�CL��̴�2�xDO��'(H��=�A�۫�dZCD�]�ؕ0��3!����N ��
��9�d^���`�� !ngJ�㈊��<� ��ѝ�A����t��F=�k�I;Ӣ*�&��ՅL�D�ѫTi�<[vo�I�w�lk\<����}4�b%� B�ϢA>�}>]>��ي໨਌z`d�f)"0����͹g-���I�:_�9=
��}���^kF%}��~�E}����CXp�п'5�@��\�(<k�n�D(h��<F����a���E�
	���|N趨%�8���& :{�A��G�o��FN���BYYd�^,>ܑL�j�w-� �VV�uacy��|/Lb���3!�95��4Z���>�������,o �kK�8���$�vS��a�9<U�����ĉ#&�����*�o���TE�QU���(��{�pGV�돇bm�*,%wg�ʛϚ�������M�]�"��O3�{�TUZ�����i��n_"�֭�a��$px8�O��]-�.���3��C���\�N	�����w�}(��^������x���&=��5Bp4<��ic�!a�#�]S�Z*4t�L�Ƭ+���kJ�xf��­�@��Y7�o�����iQHb�~�%t�M&�Ĉt&�܁�LD�}��>Nm�p���ަ�����Z@�I\���׬r��ol�>�l5|�_�D����^�|>���Ϥ��P�K6:<�>XTF�ȶ��蠖i��W�M��r%l�����]� |�wV�߈����Wb?��35�&���.�7�7n�~�S���de���
��_��If��i?z�p�R��~1h}?��T�`���TO.ع=������W<Zh?d�7��s�)�����k+������dfߛDf���d�h�8��
�zZ����u7i1���/�F��c��v;�Ҟ�b�/k� g���[��xK���b��L$���MwX�1�#>��ZZ*��cb	%�'v�)l/ ������B�\�� 4���i�0KÖ�K���V=9*>��ox��6C�.�$-F��E�h>�M֚�%����	��#=ާ�F����P����{&��-:RcDSρ䕼Z�K���XK�`.�n{TU�w���p��^Auo�eCC��5�,b-�q�?GGN�̴��:�n�~���� /�Z���p7����'��8R����(Bt�=��m:��-��8G�(c~��ΧP��+3Ϻ�'�1.���ބ�'��=d4���!��sTܶ�q@���NsJ�/ο��g^.������(� �49pQ�>l@Eb�n�;�O�GT�bw�n��2VѸ�ʤ�K݅��큄=�{�p�����.aъV���d�`�4��0 �j������N�Z��~�pʃ;иZ�nv>����_��' � s�:����� ��y99m�=n�1'�"5S�ܓ��k,��k�h�������}t=Gg5����\�ݔH�}��ڥ���C�Ҕ��*�5w[J�~��n�����v�^����S=�0�'�����dA�Yh���^�i�� ��M�2�M�隋�y��g����U��l+��V�$v�^���*b��5�~�Z�7̻��a��~�ޅ�|X�i�j�>3�����Ȓ�冧{r��ε�&��#$�`�A��s𨜐�!H�T:�uRv�RnU�LPS�]�"�=�PqH�Q�,�Š�7p�M�:�W*\���P #o���Ѱsd�o�!����N^��h������Oȇy�/4���Qe�qp�(��Vo:�d���oH���&[�����U������W���c�LU��Fm�혟8=��(��;o�5�	j2�ʩ�{1��~{)�l6g~E*���C�������K�9u����f�&��mmU׀��{F3�n�"M�$vVZ��! ����=�|+�n�O��Ζ*-�U`���`����j%�$]O�{��r�R�$m�EORC����|$p�Jw�����ɞ*������ZC��D���m�Js�֗��Nm�j�>����äT�	H���Bp$S|��+�VZ�Qx�BI4�ɶ�AHX���*�^�7Q%O�Ы��͙<y6���*����i�յ:f��^<����z��0a���P�īU@;��O]���ҍ����������M;_��-���s �؝�>�'��U�=a�S!)��Dr�`Ee��c��qg��!�ى�x#}��E�#�Q�g��:��&�w�>/�}���W r�U�����s���>F����w��O�m[��]%|����k�A5>R$7dmm5��o��� �`d�ut:1p�JNM'��c;x4��1n�6s����vG�ٯ��9�d4Pw����಍�9���uO=��+�.���?�?�&��z��&�Sw������">qh�}RRd]�IsJ�e�*�PQ�k����e����Q��ܑ�ͫ��嶽u��/N4�Y�f>I����]�'��3FsF�4([M�އY΋�����ʂz�rrڑKkkT�:%Q�;^ȫ�d����؆��ѣ�a�U�l�O�8:��𶢚��S���r�5�Н`K�p�Z\�NE�=��PG��w�D�2�I�nfb���vp����p43���Zެ����&���oM�Y�v?^����d`��h�g���/���(U�nU#�:�O�[�+8al�&�����׫�M8�������ƞ��/T�m�� b�]���'��o;Ѷ�	���-Z��D���S+e#_><�t���u¢J�6#/p�zV(8Y7+~�oS4��}��]Vu�3�d̵)�VTTx���v�������j:��Od�V�;ۛ��!��n Q��.f�uߓ���}��}��Ķm��5Bz:��̲��L����rh�!�:����"R�O9E8\��t$2�~ Ҹ2��Ϳn	���ZG��7�����b�:rX�G��PJ��!	��;ã�oQ��g�z��]�* �?�&��%L}+y����[�w�D�u(�Rϭ��z;�L/�o|6�`xhb1g�\�|5l��|��}��ݶ6䤼(� $������^����v?M�3��Dv�+��g�����g#��%W<�� PK   7��X+���  D�  /   images/5cebb09a-e86f-4cb2-800e-22da09d26481.png�yTSW7k+u Z�	�5�����dK+�т*�"�2$�!L�
���QF��bŀ"�@ ��IH��D÷Ͻqx�����w��ֳl�9g����>7湴��Dz��EA���k�6�������o��*���>?���=�'|^H�{؇@��A��W{j�<\s�W۳6d׳�c�.*��v������E���/�_K l �~�i�����n?=~�d��y�>����g{�.߱�k?����n��������k=.����yAʶ�S?7/ot�Qi�y�u�̿�]1�����_y�͜�~��z;f��ln��	�	��To��*���w�y{YJ��|���\�wr�k�0�g��2)��@�0��P7`2E��]��Su����\�64��b�BU�c�C�qs7E
{�U����|�
d� d��\�դ<M>��ᖼ# ,��m���/;K�5������k*�pnyv����ßM�GV�m�o����߆�6����m��m�����	�(e֚�ܩ�wW�^d�����RX6�,H$}� �o�h��x���X��p͎�Q���cNKCnBI�q�=qHi�e�{O�1=
x�k��U���m�n�$[G��3(��S����(WX�}�O��	��@p�9r_�6���9m|!�X!?��5>B?k��9���<W{���z��˿`��o�_� �ix�2������{�7��k��{����W��r����BE�z���V���7/��e:�I�ېc��2�?�)N�oL	G

�������/�O����"���<�Ot�"�<��,�z瓂]ǿ�ϡ.K��l�V)�8K>/��i|bH�	��w���*���w\ &�[��F��Ld��4�2��f@O���Ӛ�h^�d�+��K�������	(��S�|M��;) ������F�gAB2/	?��{��8y��v�BX�-���"]CY�����i{�\���D�=��j0���f�/q��!������M�u��>��)I�d��dK�nɁ_����Xދ�9s-0`�R�c8�@@�5����5�/$P�]�ر� �tZ�J�+R*9��|@\��5��v?��>���:��:���$2����Lb�z\G9��~\��.'�ny��!��-�q1Ș|B���_]$���	������|oS X&p�mW�c��~�?���{@�9�(���uX�MH�-�0P
����`����$/�������1��1F ����7r)D�v�s��Z|;�\h�D,1W8���gƚ���8f|��J���W���~!Řn�ŵu<��K|���ޔN�]�.�v-��r��7mrue�'q��L)R��+��¥�����z��ϑ�g҄DM�f*�r�Trܒ"S�+�#�+����ϝ��f!(7@?���9�#�?�}�+�a��כ�+��EL��\��&�I��}����I��]��g\B��Xe������)=PI�Bc��<�p��Kb�DB|~_��[$� �Q��=��g�����I2�uC����,�=0�����霫�3h�����tG��n��!�Y�^�&��~��"}d�}vxf�=<���:�G� 1��3���`�}n�ϴu+/?_��nF�޵��D��x9��k��K�n�i��+�0qa��1�y�8��h5Wb�م$59��C4����.��9��ӀT'ɛ�<�T�/�'6����~�򼚄��)�YT�\�	���)���/(�Ye�� ~��J]��*����-M��3H1�nlش-�{	0�`{7i�$�d陼'��K��R����ԣ�����]�QG��P.N���2��;��/��~%�mRN?f��
���<�WE�s-t 
��v�Q�`��m���4@FfUyrv?�m�))������-�����2.nxJ�Ǟ��߀^OJ���X4F�M 
�m%	maz��k�j���O��� l��fI_6.;�G)E=ΫM���/N���쳰,F�Z �z؅�n��?؁��< ��S���¤�h��Ge l4������,�nY)����i���8���>c�7����x&|Ό~LNߖU\��*��9.�S��(�5����^����@�Wǯ�*�Pq��R��ySL
����oâ�z�T@�� �ǯk�.�)�kD�G�e4o�����o���UT%+?5�DO�/�pƁ4����}��"�sS�b,�B5�/X�ٛ@Gr��!y�6��ē�M8�7�I U��� ��[Z��B+j��t�|�2s��R��I����;v���Eʢ:d��ЙT��ob���l�}/!�0�_P�u�[��gߊ2Fu�܂Y��.�T�����f�>�g�?�nY�������g��Q���D��R}=ax(�^~��?06����G/�v����p}�37���o�����s�"e��X�����z�l��cZ/�)<�u,D�Sܮ�E$ �CWL��U{��� DC/@���PcA3��$Z��{7�(����a�]*'��� ��̛FP	�g�G��S]D#=�
}V��.=�칵oL�\gɤ��Ìl2ܚ��N���i��6@KI��7U�>W��ʷ=�i]����Y�ݓM��[�{���ީ˕�ח�>H�=/@��kg��4�|*πTYU/n2
9��֕��^H����.̥OL��&�I���{����]��Ш��k�y[���X���d*���D؆-.*��}�l�U� ���Q����l�e��e,?��b]D~^60V��4���Ӏa�̟�SB���py1�OT�78���-ߎ�5����Dx~ء�,>@�jeSҼ���������rt*�s�!�[ͧΊ/S�F��x2�A�G9P�GT�� ˞��@���'��F�L�W1�u�p�X��YAR[,��8'�$ 2����0��o�=�
		Z�/�dvWC�O���{���.Y�4w<Yw� �Ke[�v����˝���Y�Lw��^��5oW[����e� 5����a���r�/��Rq/��.!�kV�����#��W7�h����S��k�|�Ю���)V����<+KbP��i�,2t�=7�����,g�r�S�4�՝j؝�&���X{L��^�͝�H�����浺K��,=t����O=��`=�k�i3A��xM�t�y��W��^�����O�gﱦ&��~M�pG�3a��f@3H��qo�[΁���ﾡOm%�Z���53�9o�,E�aXĿ/����Bx�_f��;>�B6����M-'�x(���];��k6*3�y��"�ץպ^��r��r8e:��M��%��G�F��E�Yӯ&گ����/�Uk�_祻����}I��hi���2o��6�^��_7U0���p�<��%�?LD����л����g(������ ~O�./o?r�}��y�3��Z:V	B6��U��3A�u��ʨd�jD���\�Κ����ӓGv��n$�[�l�} Ȉ��H�H�m�O[ó�3MI�n�Y~X�������F�A�	5�h*���U�k*�B+�7�Ŕ�(����YY�ɩL8d*Æ9ߦ}Z0A�O���N�'���r���Y9S��wnC+q�������2�>��N��R�5y{!wK��(��x�Ӏut6�^�d�_&őo;S�M�wQ���}傘ۗ�v��?�����=�2�ϛ�J2A<�#��nV�x�[��� ���]�9�]��z���,�:���Llʖ;��� T��3&�_����^T����2ET��q��N����9}�O$�[��v� �͕�,Q�̶?��܂�Qp.��8��uE�B�%5�X��nb�W��j���MY�"���U?~ j'�rA����p��&�7��,�0�Χ�K�P��sE~�*�ơ��r����ͬ�?�Q�i7��̏��:8�H�2�9/l�(H<����^��#�$;�G�z\���,��t��իޗTV5���^���l���|ϝ1����v3�[�9+�je�ŕAc��hk��R�����'@�h���FM��m�	[�b��`��baW�a=�((��2�or'�T�9�pZ����]X��,+.ˍs@+�{e
V�K�n�J�5(�0��P�$K�Գ4z�����wK��nO,!,�N����k��SE�j_��ƞ����z20�kT�l�3������}�{���R�A/=&n�b}�k���8����f��YŎ��DU�?��n�����䐻~ؘR� �j�[e4�;:�ye$"�C�w(R�3�o��9���{���=��:�6"��x��
k3������Ṗ�ɑ#p���ͫ���?12�^m���'t��2A�f1��Rf�M��h�	�D�:[�����h�:���p��>E�JuY�p�*Cʇ��;�`JLz�4�e:2������˗Fb<�f��+��J�W�UG%'����j�����Âq�l�_�τt��@ς4�A�5��|߄�v����61��Ϲ+7�[�,���Ώ.�����}5XA�)�X���ޖ��4TMWу��d�2?3.� j�!�9���~+n���rM�MG�#Z$/�¢	cd��6�}�d	��ȟSd:1��l3fN� �d*O�B�f�sC��g��<�}�=�����^��Ct���]�'��$d'�IcZ�3�ӧ鑓��nر��؊@*��i�5YyrJ.]�2$��1?��WJ6��C�xoz�qxO��-^�˭^>���U��d2�!��ݿ��5�i�իF�'��:�fBWE�撈����s#6s��:!�Xh���R�!4o����I�g��5���޾oW��"�����(>��F��=,O&��
�ݱ9��4(�t6���8��kO��}��l�뚖���B�T�@�I�|�>}d*�HUd9*�9�p�ԂE����7�^>�z�u��m7�7��;8��ksD��%����B�Cy�90�0ϲd<ռ�X��A�3�v>{��1�aEw$=�%&�S�o�:mW�b�:zs�LNc��j+����c��e��O@H�Xi�8��c� �W�$g�9�#����1÷o��&r�A�.��j��=g��MV�tSjy����ѼC�F�/�b�Q�W�@��Gy�"�Vrzώ��Y���*�6]#V�a�G���nP�^熯fl�(ǻ %��!`K�����"�{jd�Zw�8��xr�����
,����?�ԓho�F�rwc�4�c��Lb+��F�P0�[��2�P������M�����>z��|�N)OJ�eM����7�E!v�6�S�̕�#�;�/�q��쌺��}��Y�v,p�W�d�R��F��x�_�V8+Qm�WD��>X�*�wI��R��\ϭ�}𺎌c�Mu��2��c���n�L�;�������HQ�Ik�mS������ғ��*O������:���d�oE� �OǷ��'?�gd2��[�^���3�*i��lk�G���F�҃S�\�G�L��&�ۻ��u) v��h��f��+�T�����o�"F�_�ʤO�	AP�v����<�9:�wk���K�=�X���@�ުN��{��`X+JP5���ϳ���F�9?�U��a�4�R��m���f2P��Aek�0]�"z?�8��044����t��s���93�}��'bz��!NB��[e�zN���X��7"߂NaY�I*�Vj�c��i38������0�ct*���4��s�J��a�ݮsq��'��}�3���vO����C�BJH�LIP1�*OO��ARt�oc�յg&��X�EO��}����%C��dD�Xi�ዪI�|�lK�ڷg�sĺW�1���S,�xk ,X���,c�ޥŦ�c��K��=����a�}���4Y�v���T��2>��7�KX�iD�
NV��ED��02S#u=�*���Ao5���� :9�/t�����u������}K/��5��y���U�L�mt�>�K�5��'ℸ�N4'3uYc�d�г��H�rAv����9G�0�
y6�he���:��l�Z���?l�\��1�R�a'õ�(�������-WD8��̅�8p�s����dQ��-���G(����5o�����Qf��]n�"��p�7q��:g�H���?YK4i���]�4dQ�ץ��U1<��;�G@�d�x�_�6_M���'�V���r�e�����_���#_,�i���5�N��YGWR��?�O�ׁIVeW�9F�s�<mo�#\���&e��p�W�^���ź8�5��כ���CR+$���k��y��nWx�p��S�i�����7n���A�g�X�{���g��5j�����C��	")x���H$���[+%됐M����i]�%�q�j�>iꭠsނ�<��HV��OY�f�#$d,H�} On���Y��� ;g����U�ae�,�A�"�I��՝���"��ꉋD^�6�;�_zeF*��r� ���P�9�{��� L�F�$�h	�G�N/VH������%��I�^A� ь3>%9���^�;��&D(O^Ȓ�����x�,%iis�������?�elb�5Z`�]]u�[�k�N4�YwR�I�k6�Yp�C�%����$"i�u�����G��?��ҷ[lւW|���. ����Y)G�6�w�/��>�b��5�1�k��IY�#�svA3��~3��5�'�3@�_�e��!�G����iI/�d�O�
�w���j5�	�~�����'B��:�g�gB�;�u+��+Wʽ����T��%����ol�q{!~n�E=Jv���(��۽tٗk�:Bo�^�~o�*"�mL�W ���l������z�0_��ܻC�̛!z�sn��iV�C$3�Q��!f�+ -�ˁ[�d�Y���|�FS����7�����Ր�>��vv[(�l��A)ØL*�]�������&��xRnC�"]N8�N#F/�;���d�,x�B��M��Mi����M5w���(�p����ղnR�뒧U�+yD���::|,Zv.�h�ic6ȱ��v/�(��z]7�����F�F�}N�U����A=ą�Xaӝ�J6������=d\�����-��W���x�]�A.�-�1��p��Fr��-n�0Hb�Ͻ���e=��XԀ�|+&+ł{84�<�6�Q>�#`�m�3g��l���G!�Q�U?�e]o��{���@��a�+�e�p�)	�L��ҋb�1c���0�<�'���=�I��뾥����;����^��U�ǖ@��U��О�,'q���k��t�J� � 6���r�v��6 �O�&�+lm� �lTvqb.�s���|�<�����"+�Y'���>�W\�o@��0Cu�[�d1����<������q0b�����-��?��Ϗ�E���
�W_���ui��(܅��"��]�n��
��Ћ(&�/5U}� ���?��Z�?��̙.jP7J�}3�x�ţ�طKlA��m6�9ѼK��d+��6l:k/��hE67ѝ�����QY+��6ő�_��MK��_e�_��Q���j,����+i��<"@>���P��R�t?<wφ��L|UkV�	Q�Fу$^# w沼]���CJ]�Qy�U�U�	�Tͱ�>f�=���J_���~�e�m����Q(��Л��å*#d�)�e��8q�7��[lϕV����b\���%�s �"���/�:L���B�ܣǏߓ��:xj��>��_�?���Ri2�W�&�|�֖<\H)0FGy*#p;�xq��TE?fj��$"�����#
L��|�et��4�
E�zص�f���;k�ʦ��yy@�a�����"��X��y6���	�,:9������̼��h^|83C*���'
Qc�˝ԃ<�S��W�Tp�d89JL���#sޯ�C��Y�G�_���C�Å{'���!g���Wa>PӒ[!7�Τk[�s��	Ǆ31ѣ�%� r�4"֖�%P}3�4wo�@!OzSn�t�?jۦ"��!`�U;�Hٺ,�r3'���y��6���k*�Ȑ����� �N�����o��*?��V�K����&���"2�>=2������x�ꂝ�:�'����T:Q���{�i�s���;!*�ź���2;;a�E�>8���tV(y���S�#�v�N-�Z�:�7O� ���E��I,�ԆUN>5��n�U�١��F�w�����s��Q�����'|�r��l 9\�=�]y�5�c=�YsK$�N��0��݋���ħkn���B"y�77W��ߘF��2
�,i�5ֆ�*���Z�*�<߄��0}�Rcc<=S��M_�c�y��U$�e��v�}�����4,�ϻ�ɒ�pB��c�u��+ƶcw�̀]oKQ��ȱOUQ��d�Б�/�5O�N��O�.V��ѯ���簯28�Ra�Lb��ֽ���W�d�*#2��+{�+h��u��g�!y#��;����h�#�Q̖4<׌
F.z-we�>�]D�)j[,2a�0S,�����"�8��������)t�;����8�	�J�ؤ'�{���84��{��4�X�:u}����@�7�`U�2[�7F/��/��,|�M缀�F"uK���x�Q���� @0�Ǭ���2K9��Tj*���V�{R�!�X���Y��{Fr�}������҂9��z����*m��'V�u&O���07C��`n3|Q�JOQI��L%�᧥t�~�H*`��Ah��~'�߃`0���Eu�Ƨ1��v��B�y�l� ���v������Ij��&���:��V �AV�D�P�Kb�2��z�"9$�����#�l����T����EZt��n�:�O�0h�W���\}!�W��*�mXA��@r�0������߻���,B߳��G��P��\�U��_���ܝQ�p���Q(�LuF�1];��'��WEK��M�u��� �o�Zՠ`��=tt�&-�o��w�k�b>��ԜPQ"�V��N����gY{��֧ؔ
ȧ�ﭜ��%�y�5�LNe޻Lbx�M����V��qs�������Ѯ�۫,�Xюcok�$/�����'s��3T�R��Nx��Z��<2w��һe4��G�᨜����JWE�z&o���ס������<u�-g~�S�w�D	�����'	(�Mb�2np8�x�v��@|fO��NM8�'�9�Ei����u�f�\u.���u����M�c0L��3���\�\��aw*��~&5�`��`&�X}Q�@��)�ܰ=�J�m�b/�-?�f$Ɇ�є�SYVg��5�V�Ƨ����	�����T��W���ط��9�^K��\����7q�L��TqWS�0�9��]��6��~f���/���t�"":��.I"�dl�[�J$��pd����q�b;��[O���&Z<׭���&���\�L<�\�>@ՓG��O�mﮬ,��7���Ń�r��L�mFb�X��n�+�L}:�e5��7]�]k��u��;��������78��M��A��(�~0������M\��׎WaZ��?�k�C����%�S�������j�\� �e.�A�ͷ�KN�^_�?�0�l,ۊ���?4l��;��s�������c�!ǖ>������W���46�d%%���6F�M�?�=�&��GJ��{�%���m� oY�+u��%�2���ލB���O��1/�,B~�8>V�ܡ�kVZ����y�I�jnk����!�Wu���Ti�l��nz��Z��UUAe|���T�iw1�����ޞ�&��G���@�W0OltUb^Pc�0�;̺���:#kC���ix�f@��&�um��1H��������$� `�&'CrP����	����4QPn��14;�1�<��w�;'�e�=�`��y-�����-�o7#� �\�r�i��b�� I��b����eD�W5��;9�s�����EF�GM�� ����#� �苩F���w�\%�����.�5	y-����l��i�B�(�YQ�� ;�c�����l�bu�ȿݾ��Ǯ���t׼W�s[o�m�J
���G�6��Z*���EZ�BάS�%%	N("�}gN���iCEW����J�O�c6��iK ��E-�����|�P?�H�%�$_ѺoH�w!w_�R5�!s�'��M�:�&��`�D���VG8�$��{ �'����B���W�.m��x��&�T�3�I��)�ÊHg�;>X��/�M�
��7���Wj�[����AE���`}�${���DG �����]��j,E"�����}:�R��ԡM8��w;X#������]�g�Jb%�:dٺ	E��� �V�e-������M����z�����WM"zl0�$����V(�~��!S-f"e]�q��Asl �}R'łO08ZJ1ʣ
���^�h�����!�*���#�s�-��R�o�껡O��1��BS`��i�Z7\W�,�h�(z;Y�/(B�V����D����~��O��^�C����Jt��H��`��^�UZ�����A�vrHE��:��*�Zl��=F��] ��r97
�{(��80�U����׬���2+UQ�,(�dGlpn��Q�^k��V����7�)���B��Ƭ}��0�I��L_qBṄӃ0�!]���Q��<��)c4J�\D�ښY��
�]��{��&P~vR?�u�hf�/gw�>��6��e��i,y����O$�����?�6��Hx���7�۵�ՇYf�(;�Ʊkrb	��3І=��Ё���
�1�f�s�N�+y9nͬ=��jTTEh9gNs�:��Y�>��n /�rQ�`��ͺ�86Q�m�O��F(��,�abS֑��W����Z�2;�@�M��B�oL��WP�s���HkH��Ԙ/��]�;�)F��DA��w���ς4�R����>J���8I%vU�\��tY^���������T6=:@�貊<��ޤoD
�Q梲����=��\������Xw�n��yb��{��[S��X	��<Z.�-Uk
��h!�4Zχ3y�Fo��q�㎠G�[3�#���+m����r��g���5)��eu[���׍�O�{��˄��ǭk�H$N����=�h���SA�p���x,,���'�;�S��o�mIɕ8� ����^��I"*�
~�#��`�7�K(���Y�*AD���sީ:����B�Z0�K����~w�~w�� Ф2��{g;N���i>�g`Mm��d�~�������W�޹K��2n�Qb3<����687��v!�Ȋ�nǤ��(����@�W`ʸ6���ŕjl3��U�����W���q�*(+z�C���^�I)1��iQ�,��9S�����7����?�6�iJ�L&���l.���J ��IjB]��Õ��,�0q�4�ĭ�3�.-��������ae
DX���$�-ޔ����^��&���Bsu?�Wʦ˂�a�ll��Z��vL�i����}��J|,���?,;UA��DW���^%E/���/ l [Z(��h~d�=7��1�zN;%���u^KR����>�;d&�S�UVi-���xlJBW��S.�1��NUR�s��9�'Z�C�F���$��O��M�$��V!�jeEH��9��VHܲ�%E���[2�nR�ʈ�w��	@4b�����a�>�n�hY1�$y[�>�����V��$�!�$QBv�2�2A�rkT	�!	��Zx�v��W��W�f٤{O��l�,��������M{�X��z��T=������f,�}��Vc�/]Tb���	"��O6.���nv�4v�93��m�H����O;�7(MBR�u��?2҆+�w9��`���x��T����z���n�bk��m���}����v��`�}km�+�HP��ڵ��mbW,�ųQK����VΤdطC�~�1�й�z�u��2��#u|p��c�E
�L�9@磝_m��!2씵�s�7ǒŋWA���n�qw#��,x?����t�N�}�TF�pi������A��U��ʳ�74s��g��o�	R�D��R��]+
�3�}v�vG�.�KRTl���D�:77{��)�w�<~��j]Z.Ҋݚ0�t���^�^�"zd����	�������k��F0UdY1Ɇ~�>���p�|�b���R�goRv�R��R�h^$˗2��6�ȳ��RQ�س2�L�0�_��l�*��|tW��E#�S�ÞX�:����#�!ǆF��Vwl��&��[��uqd�x��kU�Rk�m��1�W`�ˊ��eww�E${`&隧/��	+zm��${Qa��A��qTζ�߿��Д9��*9����'gH�_��@���>����"Tb��E �U��܇�J������#M���D�3f�3$�y):�O�qh"F�lo�5�(�� �{wD�PK;q��7fN�@{���h��첏ަx�TO�&�So�;��_�����[�L&aP_ҰP$���{��p�E�fr<Eg�x�VT���]l��D�����V�z4;��pi�bѲO������dβ^�w��{�hrm�(e˧^�ٻ�r���B�7S�~Is�I�fό����{oH�ʵ0[���?4(y Z�b~��m].ت*�"|�����C74]��Sf�ZB��Ѡ��j���w�7Hϑ�`	���=�7���e�
*-�H�l�l�P��}|��|��ݽ�c4w���]�e�e��3V	�S�d��������������U�gz�w�o����S�ߕ�C"��?m_~�F(3FlF�9��{��Bf#��� 7�_D]]�km�/N� ��G�����5Kn$�M??X��,m�h���ǆ�#LQ�T"��$2u%��W��E�¼3;��%���O�>�}�]��Q��k��rU�w�~�ݿԠ#�Cm�&�΀�gb�B�N�ޤ;�����
����+9��)�T]:��pt?	E�q؈?]l؋?�!��y�/ߛ0TT�c/���^9
�����R�5�n�ry1Mcǩr�z~,>��u�(7@���.���>>�.�>dﻁ�s�A��ό������;GN7�I���x���(����f�0|�Z����6��tP�d+�9��޼��`1"���_t�[���	N��-�a�ￗ�?*��i!At7< �_���C��"#����6�(��Ձa�o��,K�#�b�_� �s�P���&^ V���� J�R�8�?.��n_�D�
D���h[����{�W���[���h�J�*��Կ��9x��P>��-\��rMΨg�,�~�g�$^YG�@���4d�(�g:�@��O2���8S� ߳���ë��9]�L�=��C�Ps�>%#���w�h�VV�$��p���ҏ���ύ�����[:E�g�A��qf�f���}���ݧB��� b�@t��;2�b����m�'���e��Vf����C/e�S<���B�p��`����'�ϋT]����i�y���+J��X=�:1�������6LG�?+��ڗ7���p�QL=�|�-�6~�Sa�}����?h��qh,[���T�S�QW���Pg��|~�'�ʣ�J�������q�M�I�c����L/�]y��������ǣ�K�ZxIk���'/�����'�g������ߔX_��&Z�Mkwu�i9�;s�JMG�K��3�{}&�EcZ�˃��	󗲏��v=Z?X3���x�7�o	B~����d����fvK�o�*���n[��R����29�4����df6�hl���r�14����	����'�(�L�sm��:�&�l��it������k����v�W.�|�,1:@�y󻚊�[hY/ð:}�k�m�ua�r�ע�\Ӽ�O,]xb>KM�͸ߘ>�qg��4��aW�;S��nq����ܾ��6��D�H�Tu��F�*�_��sA|��N�o�.��.�!!��;��LrI��� ���q�B��ɺ ���<u�D��<ǘ����"_
~`�>�'"H˭c�e�$G�W�0)�Ȭ�������<Öz�u�����Cu3мΰ1�Ÿn��5���笍���Ź�h���w�\s<�v��C���_(�]1!3�U����nv���=~�����b,EU�
�cDg�
cIP��"���<�Z�Yu����½JN*7���|�$�Pr��1N�����\, ���^������4X�ZO[k\7~����cT��|��{n"4�v�I�'�'�����ĉpn0e��y���XP����x>��Q���qi�/Ђ����d�Uv��k!�_I�kj�?���)xH7_¹S\ëU��`��\�p����#/�Eg��n1X��3�e�ck��ԉ��f�gic6��.ٟ2݉�����]����7�(k+���S�l�fΐ��f���s�N����	gh.�c��޸h/�B��v�s��WBw|ǾU���Sx�h,%j�^��~g��Ժ�`ڃaRlͅ2��;D}p��������ɡ���>��.�,F�v�)�K�i�b�%|��Q�2e�f��	�z���1�������r�DO�@��.Ɲ�Q�/����⿭	��}x��nni���lY�*N�	����]4�pt.e��3�/!���(V/��n:�R��X����1�K�����#����B,G��d�`MP����4CO�E��C�
����J�6D��&�{7�������pc���4v�(%���+�Ldx
��^	f��,V&�^�{ɸ����ע+'8.�f�ܤ;K �~�Wf�}�W�g/4�;KQ���[�RH� o����<�>��c��H���u����o�d߳C������N]A�P3#�D���'�A찌�������W����]����Pa=_hh4nf���I�`�Zh�ë�+������nC�>+�н�?U��C���N"c��JpZ�5u0�Ĉ�(�1���+�*Wxx�g�׽�A�Y�Ln���K��K�N�i����`��^rd,V��[%��ĕ	�串>��p���)8>5��~-��`�[��_(R!�!Y�G�j��.�
�������&lдzq�P�������H&�zЕ�l*��o�V���B�W��@����W? i�D�ME�A���*���9����T��U���u�ش<�B�	��'��hT���tV��%m�0w� U�� n�	�²��:lΰ6��}�>��Jc��P-�趁ƓPQ��j��24;<�쿁����Y�uN� �6�n2L|��c�Ze�������OyJ�I���u"�c�N�aϸ��W���
�,�(�Qe��9�_=�7�����X�	9��������r��w��o���R����)�ܥ@x�z���J̐uxn���>�&�«��_���Q���)�T_'�����,d��sDK>����zv�ܛ�n��s�!ӱ���V�Pgr�����b���\1u���*������E)�A������ȹ�öZ�v�
�wc~�����x�jpY����G��]Y��5ٓ���=�dӒ��#A�_�gWʻ����p�\�=�~��[�B��xZ_#��\;�局T� 𭀓�mr����;��"w3Ȇ�&����G�{�Κ��vS6�=��!�D4�uY��8ס�/8
�Bk�ˀ�"i�C�e}��M1z73A|Mf��ҰY�z�@y��nc��~�¶� �ڟe�o��<s�|Cs*����r���"�۷^tS����3����&
��P�p��DHA�yj�'��W�َ�/��
R#S�F�t��b�MP�L�Ȭ����?�ݑM�%�>��B�-�����~�:��Y��CFݺ�'�FH��m/���&]�cK w�4L�������c ��:��� ����ox��� �c�l!#�}��χ{�<5YPk���
�&tU�������.*�O��*���0�����G2M��IPd���H��@g
�BJ�'V������d.��o$��=�V�H�{��9��--~���5��p�s<��OA��	�%=7�T����T�Q�v}v̄`"����i����.z�����UiJ�w��(«���q��� �a��]�*#+�Q-��Q���uZ��� m{�ؐ߉qة�i�������:(�*x�j�b�|&��;�_b �����豙9�R�����qx�a;a�추}����s=�{����x���4>��&�G�I����(t���v��$���?�J<A{춤�7��7��YH{��.HQ��y���O��_��قt�������6��%D���1��'E�	���]�
S���܃߹��?�Ci>4W�Cw���rg^��xڣ�v3P�*��LD3����������{>S�Z�ڙnX]��xb��s��Q�V�R	���a)�-�[y\����B��뒔�^��i�ِ=H��PX�
֣���/�|y�L0��#�h�ɁkWf��<�Fח(��SRj%�|�yø6��w���hc��=7����Z�Z��/���.|����Ԃp�-mݝ���:0=I (��D���5�Ѝ���#�Z&~x��_��)��`p`��&(Niݧ����w4��ܲ�o=��9�����TBͧ��o��_�� �Ss>�Z)&�+�Q��f@��VN|��i�a�D���w�A�~*�-%���f�q��] �㷂�uSw��2�ED�+���Rv4#���y�VD����s �`wu��Ai��ϱ�x�8^Tkx�B��&�=rө6Y�hH�P�F�YG�U�$�Z)����ۍ�.��gO����.��ʼϠ�5�7�͖2R�����k����n����?���T��=��h[]@�ր<68<5�y0���H}�a�ƿ6ȱf�����z���_����y�\c� ��:(�2r���/$�Vx0#���Y��ꚴȹ��� �:��q��\%,�|*%��.�_�S"5�����1�K�f����� ab�z�U�w|*�� �G8�u>+�?G�]�Х6H�)��/$H��hOp��tZT��Xj��Q�OQ�rȭ����z�~ss�|E&YF�m��}�R@)�3`�+��F��C���@�A���x�J������o��؉q��5��U�.A�,���O�8�����kL����u��tR�f�C�9�K����Y5Q��f��L�kf��%��,HF���'j?��(�+����JI{�����A^̪�:����>��'�E���Բ�SÉK�s������0���H�6ۏ7�/����=�~W*{�>�B�;z*�?5��zq�v���$UR����BZ�d*�S�(�E;���=�OL�`^�ߧ'%��A|[�V��‶��O�/��������>>h|�s�]3w�i�o�\9:m�&y*g�TПL��ܠа�4�M�v��&��lt�;��XP��f�a�j������t���X�r|$_�XR�3��y�A	~�k��I�˚��g�g0}���ᆪ>�ϝf��#��h���1�4�[9��.�,���c.q=�cQiD�"�:pݹ�Sr��u�6�3���n pD��DE��8)6rt����'�p5N���ظWt��ҹw�?A�6��ā=-�#��V[�>1Y��q�󠎼�Â����B�u����v�-�3��
I�r�Ӯ��[��*��F��#���@�~�x�P��R�/T�d�����10�=?�� �R�ٓ����I96.-271qH�.�vJ`·v&?��{�s2�����ʘ;XW��JR
���L�Qv1�>~8�B��\�9Z�38�Q 662��6����(.�c�\�|wV��y-��1n��8���G�e*��}b E�u}�������eϞ(�L�Cς�&�!��V�Д�tg�n���lĳ���,�EJ�YJ��v��J.���v�ƒzD�����P�q��<�w�|I$28gBf�o m�[���פ]f�P��l��ar�n�ׯ��-���ySnG������M�y5Z�xGZ]-�dP
<s��a��B������tZ�ݙ�w��x;�G��T;�R�`�dW�˧�ܮU�O�8T��i6���ߕ�)R���E��(ʺ�&�>����o�
��A̭�X%� �uϩ�<�)�Y���a��U��L
��a�:l7Q��Ɂ�y0���T�n�0E�����\����t#������k܏7��k'��K�j.ж����?�Q��E,�B}H����&���� 7!�C���ă���]��Etg���7;�)d�ڠ�"�K~I����E	���.C�l��,��@���;�����&����K�8�]Μ39�� ���~T��?��mOj*��hYMڴ��Z����(5���ff�i���7�߱���F���e�ܷ�;>1�����\5c+�_���l��eh�4-^�O�#��R;��MM��,��8_�HߺN���!`���8j��T��N�$��� ���WAk�Y�5�H4�M�u��Ű���������Kdlԁ��R���|-i��p	����4�x�q���O+��s��Ccq�،z8��T��h��3FpP��l-Rk`bbҎ_�VϢ9���~�ف*j�h]@��i�M�����j}3i��.�L�⍸ۆʒ��g���?R����
5�F��SŴS��G��&s�%�؍��[=jHڅׂ�f�%��`��:�V�(V�"8T�s�MA#l"�X谵f�hE�W�q��*`P3Y�:vtkr����x���RvxL��������Me[�����+�s�+2
�� ""J1b(�0#�:��A��Z0�6�U�Q�9�HW1 "E�^"�`��[B@HI�PB�w�s�}�?��|���|��>k���w���0�E ��b�>���f�}�J׌Ω혢H�����"�(�=;)�B�OG��h���[�ƾLÕ�[�i�e�6��!Ơ��LX'R�����L��*���#[ ���(i�@�M�Ǔ�lI����w����*It�2���_,�_qi�������w��_˪�峁˼(�+G|4G���>�5ޠ�Z�k�뎩��ʾA�6�IO��K� ���i�چh�S#1IJG��$�3����x��;�3�f�~�;�H��o�鿁3Lr����a;'�Ľ��X/tLU�:����N���+��A<����N��j�Hc"?jo��\[d	��mp��F12<0�67q"�b�%�)y���|�&���
l�ܨ=�լAY�B��M���M�Lg�OR�tZBC�5�W_��~B<�;�ݝ���oz�����z����K��i�m`��k��ȇhّ����� �a^h§��U��g��g{����7��������vz�ޚ'|��� a"�g���`����SV�L4�Z�b;��]�m�c	(T��г��l&L͛Z��V��݃ڪ��Y���zk}��+-��L�Qj�`��Us�����=4i*�ܴk�L�U�;��HC�Q�x�4Ӹ�O�<��w��ʑ%hr���HΛM̮�>% �䛚����Ԫ��	k�k#�3Ea���O��{q�~;�Q�0�-�J/V#{u�����K�}:�+�%vh���L_e����f���;n�(�3�f�F��W�����������Zx�BWؕ���f�of�q���Ӓ�I�v/n��[%՜/�ܨU4x���R���2�gO�.�G�R�p�ގ�q��)�6 �kY����$٣��#�/b˴_�k���c�������_����HTF��F�<cN�i	��e��� &r1�Cqdۼ�5n���J���7��ՠv�k]+4�_�q�ablxX"��Z�Y�m��uL�&1y��^�r<��Uk<NtZX@��e7������ͨ`�V'����˦ui'�xy}c�s.D�#.�@��U/�g��h�$c+ҋH wt;�2�n��U6� ����|���z���楳"i���3_U�a��ZV��\�Ò��K� ����v7jxdg����L��5�@�F��U�p/Y����ƍ�S�x�4���y�7�1�}�;�7�c�t��o�ε&Id��vSb����;�ƀy����x����ܐ��dgb�a����2Ȋ�[3%��W�v*�x��-�(����o'oC�ܷf��M��N���!�ԥ�YX��")��f�w�:�e���r�pc5�#�a��������u��8R^0lQ��ޮ����>8)H5T)G7m�
5�o����3y�aQk3c���#��&�gw5*�3a��S�޾���Uʈ�a��S6;�[��ns�@U�Bgc�����EbXf�� ���jO��[|%ju{Be�W >P��p�V�G�[;/s����*)]o�>������aL[y�
����{���4�s$AK����c���g*���Ab����TI3�$���$v���.���x�Ǉq����j�"�X�&;�Z���1��=�`7}k���p�P%�=<�ȕ�{�Rn4��|L�$���gMX���h�`(P?����-���G2�{iG��R�?���/��쎥���4�z�_��~(a�%%xCh�`MIG�,�7���B��.�"^s��h�w/�[��4�e�~s�Ɩ"�>�5p���7����kヮ];A�IF��!�`��3�񺒭dT�F'Y�2>����SV��Ǐ�ێ�t+�R#�k˛ƍI�����7�xc5*(���|����ONĊ2%��%��ȿ���K�c���e�SY���rT���\�U������V����"�[_�FӱZKY�g:qhs�+P8�G�
����Qb0�5dP���2�C��Q�z����&���|�ٶ�~s��iw-Xd.���Cp�B��k�y��Wg�z����A����T��3��+F0<��E���3�=�=�"U���� �(6����d��g�>5E���t\� m���;2v���"@* ���I�1��4�	��U�?�Y�˨�G�����*@���a��%*�O!��v�U(`I� і7kh���v�T:�ٖ�g�u|k���l�\,�3c&��x[Hh+_Ur��|������������H�L?#�3�5����mc=
�o�!{���Y3�/*�GN�l���	.��=|aKC�5O�kd#]~��6h������NjD ,-F[}ܪ=*�V�I�A�Y~�]�ۡ��6Ho�@)ϊJ�e#ms����w��є�̖�ϽiM~u_�7�Q�f�C�s
Bd�G�J��̳�1 g�q�wO��湠���_}��6�\�ffY����ؾ��h�/�Xgě����E��,]ZPp�-�@�� BmF>�%c$�j����ѵ_h��dC( �}���v�(g<]��K@<HZC�]뫵uTmP��NI0#V��D�5����7�ۊLTȝ[$��ɜǀ��
iO��%�^� ��oղ�0������.��h�%�'�g�Ɗ� i���~�Y�!�k���7;��� 
 ����Av�c��
�8���N��ϺcE:���ϻ���1ό[I�K���:#i,����My��p�v���2T�Yß��o)1	A��aF�������x<�q��(kU�7D�V	� �M��:��D�^w#�0(r���O�,���j@�
��0+�����
 |��i���p��f�-�E��J��Mɍ��K0j���C��~f<csb~,��xDŤw��1%gp����gd��c���y��]P�2tg|��b���ț�� Y�S��8�<i��M�(��]��x���.� �ŌO\�w:��AO�� �?���h�2�c��w�wu�H�W��3�Tέ��{�] n���rݿ�a	�O��*�~i����|9�>B�#�La�z>>Hr�!�q�oܛj	4|�|����sv�d���#�������J�@́�����;ekm��2@Bu<FK��.إs!��E3����@~3v�~��A%�0@�G��#n�(4�k1H�*�W�Q'@G�yP,&�ghj��3 �W'y,���2����Qa�MĻ^�ѕ�d�F�����2��a0H���#�Z���}w��Q�ڋ�i���e��n����p��砀R[twl�O�xf�մ151������/����e���6��d��,��T�>,Z����{A�}�?o7L4�S����� ��u���Vgu�����z)񹒳#�
��$��Ǩ�mFM��ۨT3��1��o���r*B`�ǩ��l�9� ��!O����b[=�\;�(&v2݉^)�-</�"�e1�E\(��}����S�&O���E��)�\��m�B�  ac�u�bC����7`��Lb�)\�=#ǣ��81\W������� 3:f�Z^9�cw�[���� ������6,'8��+-��r��
��pQ>**�����
7��,�+�kw�w*/��G�K�` ��"O�Z�zP�$	cq��V���x��d`
�]����]Rfa��LE!Pt=x����Z�/��s��-CI�
n$$�B�� �h,ù>n�u���z�ºJ���	 �v"�!�~6LU��^�͊�%��Z��K_ *T=��b$/x0�0�?�>Kќ����B �M'�T`H����j�SnL��8Hl3_�>�m��7��t
;�a�AdK��}��&�z���C����r��n�Ҝ��{q$��9� �+���\|�
c��ٗ���`�^mG���<ި��"z���Y����N�%�\����>���o�!��?�pZ7�`�ô��wJjn���ܻ�9�UL�X�R��YR�_��:���Pٖ|y ��t}�i������F�xC�����q�'�C�Ca���5|�O��Z ;K<Q9^(1�����T��W��y� +3�e���t���!�1n<�W��Lu��v�!zwl˨���2�����Wq�z��F���3ޙ�� �s�,$f���+ ��(��oj����y�W�	�.��Y���#xw�Q����1�  O�C�;u��tl�(�󭻘�9�co��e�j�T��y��1�	zH5#,��ɡ0�IF|�s�͖�ɗQ^�����r���n��@����o0�j/Rf���;Zb��l�c�|vm�tc`�P\/Ā��]� ��!Ts�\�'A1�� �(�x�S�� n�ѓ�1�?�5�0z/叝�����|���a�X���d����L��f|c�z���8}��������3�ȗ0xL3^�"�m�$�c9F�=�<2
^��5D�eay�I١-�t|M���v���q�Co�z���շ_}�������_��_����o�Ҿ��+G������F���]Z�>5䁕�����__���չ&iԯ}`=O0
��J�7�w>v��|U~�0��P%�g{F�Os�xGK�D������ݮIQst�=�]lί,?�28�e�ш�F�O�v_,<�-N:�̰"5���[��^m����C��aO�۶�a���N���A�5T9rW�-϶���}�6z�®X\ά_�x�Q@uqĽ;����9����E~�3v�J�OB&�� BnYYF�h�R��r�|z	�E@��_g�i��-#?R~p�O��M��o���Z�0��@�ь� F]�	�����6��%$����~0��O��Ԩg��*��{)�1��3UF-u���»:��L��	j�iIl���~�HI�����v��K��� � <����u�L{8��W0��q>�	��a��!�'�D�#҂*��@�,O�v���9��z ?F���e�'V�
��p]֯�?G��,�\���������ǹ�'0��a�q��6�������x%0o)ݺ4��S��t�M2o)���=T�O��G�+��zĸ'˳ꍨ!!e�0�cN���Ӿ���*�J���)#�-bu�ܢ԰���O�\���T8�ed����h'c��i�>��v&��;�T�j�+�k^�����[C?�%F�/eK� C�tU�w�BdBY~����+���4�YC25~^s1�
_�T��i��1ة �efh�?9OO��z�u�%��|�?��nO8��"�ax��.U1��y#YG�ͱ�������R��XF�G/T��H�ϕ��~;�~�$�1�iL�Yܕ�u�X@�g���ZUG��eU'M��? go�o?8��t+v��E�@b���(j��ä�'�.�<Nh����3��gB]���	=�>���}���U�Y�U2������|�)����^4���{��Vo����VVgq�FvD�t��O�:�T`*�&X�G��ʱr��0��LO;U�>I k�Xl��ʕ� ���]pWb���$�ID���Iv�i�h7�C7�U�"�p6�q�w�U�S��Y��F7~�"g���4�rgUݵ1��%j����C��1�y�����9������39��@z�b���|4�Ǘ>��er�G7~��� -���<��q�9|P�kݎ��Oһ�:�{�ʮ���#���B�V��3��/SaǈbdiA�)1z�B�&ܔ��V�6�{��o�d'*���F�&�7b:0�ڦ���akW����F*<�ꋿp�j����6l��ZL����(_�3$�ߩpZ��q,?hߓ��KH^o4\��IY�n�$Ͽ�ɃG�0r ��8+ݎ��uv�?�+��o�h�\�R �_K#�N�-7���"�^��k��L鉹����e��>VР�0g���Y~�)7ZJ`�
��<K�|(����Ȗ��퓻�\�b��d$��ػ��s�m������1h� �T3�F��y��k2�,m䫹ſ8c��r�ȷ���i\��j7 Օ$���n��B�D�[0�s'oIVC�IDH���
���7n�į�ni���շА�K\Bn�E���Z���b"�8����[���[�A�/	�V��;`�U�������ḱt����'Y�b�\w�f(����1m�i&��ލ�(����!�dH몥�[~��	��[C0�*Վ��A��pȚ{7j�<x:��(HHu4'�[fP�~Lz���P0v@;"�2��G�4ǽ��цG-�~�j��F�z���.�ye%�]%�_D-�F�7_�ʸE��d̶j6]�@2*�O{lh��y�\�N�ҝ��R7Z��ep���xu��(�t��e54���@�UK�2A��1����]�	�y���o�^�*��D����9	F�Wj�Ѩ����W���Q�D��T�	��	��8)W� ���;�6�6�
0r��lK��s l�ү���`�x�Mo+��,;��,�ӊ���w��)��]��F|��]�g9�C�+k�J�8�B�jA�Va(c�^`t��>9�5'
(9_}R�|2z�tX�o�Nk�- ����ֽ��{ҧl �`u����ͬۡ.G�^�eȻ�6W����O���7Q .qK��Qi���e���b1�Ϊ�㣖A���������k��I�G��R�I��f�>�l䀉/b[�cG���b�C��O�����}c�]��B�����1y�BW��4��a��~�6';���տ�V%��EMk������pR מ��4�F}�q�v��������/]m|9��55��YD2͎��$IF��������2�Y�VB������n+�%�ro4̑2����)}u%B�"�`���a�P�����mkX�Aއ2�:o}�������@������6e�ŧ�ڻjX��Q��v��ZH�l鮗|'�Y���)79��5|�~RN�%�7����e��Q4���eTȁ�n��F)9��h���!{��^�i>��FE��&w���G���mW�u����R���қ�U�6�v̐�����7Fv cO��M�H&��+c�fA�#���~�J��T���P��ڌ��Q�<�i��1�L
?�u��A�(%��^_����$�q�z���[��&�c�`"�e{�=dp�a
"WZ���z �[H�ߞ=�O��ظN�\v?>��d��<�٩ۏ���#��N�;� �P�:�H!D{�$�Y�HT8JO���	�8�j04�Le^��E�J�<X�c�R�$���޳y5� e�sh�����you;�|��'nr+����;���q�9䭪�<��1��Z�9��a� ��>i��#\�˔��`DR3��&977j@tҫ�k#�*��fk�ֳ�s�_�Go|٫$-h\LwT�	p�yX�{By���v�M��BVw�.�k�� �������_��y=4������u���%������ߊ@�H<^5(�o�2�0��՞�)�ҋa]Y�j�u �&َ����$$�4�Ƨ��[�0	��_&��`hq�xr�M#�z���uO�(��2>=W���U��J����^�<�>B�N`�aV�����W}ѻ]n$4�GG�|.l|��8�s?f���럚eT���SO(US�,Oc����2�FƁ��@��0(��d�ضn���v���u+��B;Y�XQ��	���_��!�!������g� �)����7��<�W���P�h��(�4�<ډ��hz�F7���=�D��eKRӄ�.^&�C��򋻋N��`��矚Qg��*'���׌�1�%��*-�Z�ږ��J��'9���-�1���v���:P֨�:XY�=@CXS�xC4��d�}���1� Ð�����+ulA�Y��J��hEQ2AZYv���l�Id�䞨jF�+ǻ�!#�~)� �ƛ�<M��zK"#�X�2ΠM�t���@�ȣ�Bj*3 ͜�(��p��a�2B_�R\]j�;p&����䟠8r��1MU�?�p��m�dB��)�G0�rn��ܖ��C���C���č�v>9;���v���(�~����٪V9*vE'�D�Q��z ׁ@/4x�B�[���ض��q�@h A����{�Te'Nv�Y5�jΧw�T�A$�q��0��(ޮ�%�3�����+'���b�;n~=�q��$�Ӓ�o�v�[X;rs����E,�Ez,Y��5n����_�|�9J�܄�L��KI�ƍ��HWn�o�U��+��r<���2,!��W:��?�~�d���d�_�jF#��C�� ��B�L�cY�,h�H�������Sɘ�paK9��J�t0��Q,O����]�B����T�|�AېQ�����Sc�)&�:(�{��M��3�!�1*Ȇ�!Z�=�hD��L��gO:���X9[�kS>�Z��XZe>�l�q�l������fR
I_��Q�,N�ș�}y�h4�27>���r�Ʃ|�i�!�Uw�o
jY�@� ��,&��+J>�{)�k�j��xH��Z�ԆN�ذ=�n��!1��˛�Ι؇WJ���ُtw�_qn~�*8X^R�='OXk�0R��>��9���L5��gr�m��d��qzϩS���5Z6�_H���Ĳ�S짙�Tu�z������`BV5�}�tsD�\���Ǩ��o�+�ygl��*�+'#���x�Ǭ��{�|zW��B�ܵ�/3��No\��8�m�\��j5cD1�����f��8y��GhPE��SǗ�Aɘ�~B��͵D��B� ��޴,� 5$&��Q�����֩Ҫ�R����/'@:T�)@N�sc��Z�Sc��-���d-�𙇘0s���c�6ɼ�WS�ސ�÷��Jaȩ�"4�����~�iT������2�G�8W��}�6\�n��}���������r�����t5�Yn���6�F����V�e�VR����`��fRh:�F���1�dxEԓ�f$3yp?kN�n���@SJs�<o���@�����u ٹd��[��WԻ�Q���T�a�P�N1:�u:��t(BT�~gkO�#~����&�2:�XF��Z�Q�����s�o<qaV��#�[�{XtT�<o]��p����⩛x�'���m��<�V�C4��e
)� Ħ��h?=���K��@�$��V��]!�������W���|(@^aR@x>�����%��񫔍�����(����{Y�AW��c��@�	�7 � ���]�a2в����k��-�N�a;����T�5'o�=�9�b�f;�קE%6Fp-��$��]��^O�=kQbֿ�S�������!F�Mû?�Q}���|*���⳨��oW^�(���I�_�w�����V��OƊ����v!�ш���U�9��n+�?���õh�vj�(��=��O_em���Gj�c��/�����܊�(5�zܨ�(�����9/A
�+&�~��w����jK��B-X��Nc��:�W��?�~��"B񄳀db.yi!��coՄ�)@�bp�ċ��ikM��&`9�
�g�͑{J^�'����GG�b+b�w��b���~?�(�E�MY���͓�lm��,������������g�n��NG����^f\���<�#��'��/���J}����礶��+��
�D�,��;qP��rُ�K��'��q�f���	�����ۭ�h�,�Tk;(J�1_��>��U�:n��K���HnH�ZIn�<y�Q Ej�(\F�_�cm��x!����1H�}�n�l�w�7\��n��;��&g������C��8-�[/R�����c\-�p�>��VW�ۡ�[)�hۙ5"�<��JRc}<�R%�B�Pb�~_I��l�Ju 7���LB��4����R�#��T��<f0(I�j�z+��Oj�)�Sm\&������ 9�a;l�H��a�h"�h�l6A�1�$�G¥h�C'�Zw�1J�/Ny�^fZ�es����Wݿ{w�Ġd^��9���ݠ2(á�����;f���Z��C���D����������a%���_M6���%�}��`ղ� *��4�ί7^Q�)j�2� &C.w9���t�F_���J�:��
����k�����bEcs^B�v
5�{<��t�mii��z���?�{�+)nF�7�o�m|T�m���^�𵝴�0�XcZnbe��Q����+D1�AMh	%�
k1���{�˨Tz���rg��<�I<*��)���*g7~�x���<L*���Z�+۔�ڤfU��vSӑ"D1iŊ��;m�3~�W�ӛ!F��~�_��}�\��j=�D����{ݪh,C��蟋]�"xx��}^��#�,�?̵GCNiI��q9QF���uy	]�i��P/55q�O���}�h^U�HXr����c;y�Ս	�4�8�Sw$a>ۂ�ɻ�b@�����?�7'3���AԴ��oǊ����r�Q3>dQ���F����T������lȘ#*z��'� +�J����y���7M�0����-�X9rĠEO�+7����$�����DE'C\ifb4�բG4�w�=}nϕB���>Մ�����^�C��[9�!943
/D�6����r�$����2c"uk�6�<}fv��	
��jX"։�Z{�=lH�9/7 �|H�E�UA��U\��� UjÃW�Ki?n��P��Z�����+f��ԆxN�K����	x/2E,���|��̉�v�о�,v��6+}Fj���4�]t�s�{u�Ǝ8�+�r��`���N4�k���(4}<~=���5k�}f20tjǓ��q�]���c�dyD�N��;r��/M�L0�}?(!`>��1j?�
̉!8/�G�p:˝o��v��U�A?�3"��x�!�(�)�ۊֶ"� ��[�0eg�_���-���R9,�"p�X� ®��͍���y����oW��؏Yڲ��?��+�5���@���;��l{�R�y���8���,@��0��@B�;-��_��b(��J�'������;�����J/�ڔ�#ϻ]�}��b�͛6������~� v���Tҗv�':/ X��֭l����;��n�1P����>PX��UMj�%lK%�%��.@�H����"ۜoDxF=��a/�
����tNT9�ݺI�E�?�t[��aɬ���R.Ʊ8��s}}���k.�>`���>wdW/��M��H�̹��V㎅�4��
	�,��Qv>j�M/������e�����ix%��uy���ǎW锂
ĸN�CD��R����{�O�P��H7=/7���O>���&�֨�+*
��{�4��iQo��b9@�4'��Z|�4{�H��iv�������A�n����>i�v�Q�y��({0��t�3B`����A��x�	�G�8��N,�$ �@Zb�!F<X^�O%���ԍ̄\�>X�����W��ʬݼ���L�u�g~k�|��3�
�S1s@h�\2?����)���cU:�^yy��lA���dV�kj��<zs����x�I���,#�@'�(�f�hF����L���p�79E��k���@���?��lF��d�z�a7^�5�F�fB�n�I+R��ҭWn����z���hi�F ����
�?�D��~.�g=����}n�ԅ�fۮ�
��)�EkN�Wo:��آ��o��ȑ���Xh?�U N�XӬ,O6c�=>�&b��,=W���{�T��#E��:��5���˰�&*�jxP��:0�g��%��2�ޗ�S3"̰�\�|���#I@m�)�;F(��83#�b��Z�-�G7aLF�XV:���)��v�ތL[�<D�c7���^����<{-�-�{����S���Ճ�@�I��sxfƘP�
�2KHmf�&u2;��)C_��-���#ݶu�o��?��Kvy�=(>Ɠ�-u 傕�]Ξr�3o4��]�hL?�n�ퟕaP?�{5�Y}�9�߲v#��/����g�٫�qO��E�x%�_Ց�����B�]Uv�����t������;3|*ŏ�樑�G��9d�O/�_��ͭ_��=�LBdd�Z�k'��9�լ�\�9�ň��w@���r�c
̙����+U����IFw��K�v�v^�����
v��5t���/~p��_j\I�75���&����`�D����2:����\8� �u8M5�nB��Ix8|�Y���P�I���ثw�d�E��E:l���Ϸ^�P^�h��φl>A�[ ˛O
Pc���0�������Wڑd[���^�ɨY�K1\�����0�Hm_;*�=��Ԉ���U�v��OO��
G��ː^9�̐\w�ۮv��y�NUp&�A����Qu���Ʒ��������UB�lK�u���#=`�#4���95��e8�|3~'v'5�x_�|)� qUv}��^��qQ/��#�je��g��ވ�@����bJ�5b_�-�FS'���3$v"Gr�nq��ה�R�����xL�*!8'��v���^��A(��'M�"y�\C�k��"��RVc�,5�x��4X�[W�^�q~j�� :�=(�nG���>ܴuu�z���l!y�lH���Gi��_ /R��*���'���uU�%�4P1��T%Tu �m���Y��73&i������<��)R�2Q>[ֲ?�W�坨��4�G�S�芖8�[ci�7�=}g�</O�Y�;7�u��U��q4�鲼���33�G������vo�8��Q}��$5|0�}�:!�G���>�lg�^<64c���A�m�)Y�	od�x�U(Tй���ѥ��䫒I�Ɗ����/w*�d(�U�~��K��>�K?)-8�Xj��P����9^���YyDsc,7GwEy�+Ɲ��9��\��� O!x�0�^�����D��@F����l�o���\�̃���6O0�F4i_:^%W��n�X�#��>9�~*SG"�XƸQ��ah�Ȅ�7G=�'7�L��9)��Ș�ЦM+G�E=��ba��Y&�mΧ��I�Lo��Z������iֻ��l�!�i:��{��$;�A��G��a�H�lMZ]	~Ӎ���bk.,%ͤ��/r>^��qܕ1�=�GW��|�B�u�n��#���zEmR%Z��B\(���rN�R�����ϗ5ͩ��_=��U�� �8�'m��h=������̫#�z���Db�D��8T rb���j�K����N?![?���b��Rh4�O?o�Tdq?�h��P(�V�ԍ����ʡ}�N�w�h0b!�>�DMG�����A2�Llc�iE�[tz׈��;��\����u���"�i<*��.j�����Բx�wV~��	���5K���x�BظG�yy�2ݨE:�'jST�H�ۃȖQ�鰶b՟o�P�,f5�:���>�n�Y���~+r]=S:����!���a���������T��F��3ٍ��g,��o*::�o�3b8�+�\�͈2���'!)嘒,op�b�	�Ǖ�O6 ������.g�Pm�*h��?~�4�y�hc׬2(T�|ҀUΗEkY-� 9���?�Ċ�[�(�1^m\ Hᮭ�cVS�oZ�~�`398�A��{�v��z�#']�8���'(a��Z�f�S�P�Tw��D/���t[��kǽ�ń4(�+4rH������j$�+UU�Zb���'m����m��)E�3_!�l&�s��=A������;��'�; $}�Z�����9C ����+�@qI�=�+u[�M�.���x�2�T�L�7�D�o������¨�^?mVW٫���(���I�$d��E�w#�k0�����Z����V�T��1?������Bڰۑ�]�!���;Z��n���������oj��+U��۠_���WPai=V=�kXDz�|��!��H��3!;�"�<�*����2H�J� ��o��w��P�~�oj�R"�֭� sj�ߧ4���?B$�?��L� Q�ո�Ο
HR�~�iu�˯^b8��S���$�+k�
43�.�6am|1�6��Dy�[�Am{�*�WF`�MT\ft1��J�!�{���	�q�i���O!K]P����4�<1Z� 	(%= ��"27�%�M�"%&�S��p������s�ܑ��1B1O-��KKTk9�~���Klc���LU!̧/Y�o�퍍�P�+��Q%#ϛ�NVU�\�pG��$4���v����r.m�f�Ԕ��[�KoO�7�U=�h��8��*J�����*�F#ga;>��x��^�Ч!1W�{'8xZ��J�g��l�tzg2�14R��(!6e*�٨w�����h����Uey�����j��3.�2GПԚ�3։/XVK'ͯZ��sٛ�l�f�k��,sE3��F����٠�|{��|�[�c��
�d��y<�pr���d.����x�|X��;��GΤ6F�v�p�,X<��l�A�5��/�/0���Yo�JWV
z��8n^�}�ǜ�ңۅ�!�z>��͸sT�y^]��j�"[2I3�䤦.Cd^��{*�lvȇ�A>�0'�=�L�>G$,�'VD����pԷ~�iT��-De�^uZ��}C�k�\��QG"͘��q�{S��5��O�h�D.s�*�n�,qI�u�&�9@�PIq���S'�l�^��`=͂�B(�Ca҂���=(?raOB�}�`��WH���Ygd�%K^��X=b�]�}�^��гzT�R��D7���M��+�O^��Z�-��h�D�uܝ�P��V��iY�� �}�e|l�U�5,����B�����$+�z��aί�I���k��{f�Y#�r�a����]��d2�$K�QR}�C���Ɯ$�ht'�g��8L�����b�J{�U����KDft=71쨵e�F�"���ԥ�{�)W-ԽS����-�P�ɼ7�Z0��XX,l�癬��}e�7��5_%��28[M�^1�H��@UU��i���2 ����21>��Ȉc����fh��)	{q̯��@�~���E�rZQ��^�Ȧ�}Y��*�v�4�����%���R�#-�I/�Q:��;�lS�n;}����%�k��W.{�c�7}?n�Z�;��'�q�N��#?�����5R��{~�~m�� k�I��[py�_�O��uK}���Qj�.t�ￗ�pZ�S���-���B��/��B��/��B��������oRRߒ� ���B������S�J��
1�.����ߌ��v���p�c�OJi���no����5Z���.5Գ(_<�>�V�xO3rc��`žK���酱��^���>��b��ӧR��㗖�II]�i1�zG�(R)��MMbo������B��/��B��nΉ
&�#K��=�I!ӛM���������Fj~~��y�*�P��V�pc��=�_d��vg��#�S���ۤj?������x�tU�[vm`�z�\�h�)^�9p������K�Z��2!y�I2�g�e%s��yL2�%ɜ/>����_|!���_|!����fCOwJ}��ڴ�e���k|+�f�z������x!c�t#������w֝mj|\�,�,��������K��PK   7��X��/F��  ��  /   images/7fff522b-95d5-4303-ab4b-62aae53cf766.png ;@Ŀ�PNG

   IHDR   �  w   `�3�   	pHYs  �  ��+  �RIDATx��}��U����קd2)$@� �����T\�����b�����E,��P�� ���R$"���H�(� 	I������=��޼d2d&�̲^>a޼y����{�=�{α�o�oc�o����7������a�mlpL�X�h�2{���;��C����vuwT������M_r�G.3#�7���{r����S�ryJ:��l6���^:���4	�V%�;���+����_��W:�݇�xo��<^�̬Y�h͚5�������|�~t�Yg^~�Qx�����n�i�뮻��<����Ţy�G�iQ��8��>��J����EG}����z�U'�x�[c�[�0^xᅶK.��w/���S>t�G���_h~�c��ܹs�������2���$��r��U�VA$�ʕ+m>mg���=����}���a�4I�y�w�%�\�N8�����{  �"���ðx���Xx�]w-�߃/�˟�袋�ݒsߢ���/~����2�K�~�s睷��OAX�z�J�P:cӚ��3[M�eT��aX�:�Y�g��]�����y_Zh>��C�O���3�������y�{i�������ۿ��M��ַF�oB,�H�;�:����x͟����o^�/|�7�cKq�-B�?��>����[n���V�s�=ȶ]�
E�811�T�O�G�kS�=�����p���}��ߵ�#�M�_Yb��GWg�(֞w�9�����O[y�������%�a���i&�7����'���3�8�ܟ��'ߦ�<6;a������΃~~�y�O}����I�_���~�dSG�'�Q�t��~�_�۟�̙���t�9��KO<���7�p�?�V?�p���[�x��)8���8���E���i^s�5�~��o����1ڌc���W_�3>��;������~����W�d�!C��Ü�cvj��5Qlx�4�+Ez׻��'�x��k���eq��%�\�Cڂ�Gi�o��z���;�^���(0p�DI���QVL_��O�����f#�~`���8���{���ݱ�ڊW����5oGDF*���6zF�^W�"zz���6���S��<������k�|���?�����Rɣ�O���F+8��Htp&�f]�7,�~C�al�`�#�J柿��������AJ��S�d��XB��@N������<�0`"��R����@L����4m�1gΜ%�C�b}Bh�H��燿�c�l�6�(�_�hQ�����	��,�q�Y�����6�=���a%�f�����,�u(m��^k4�H��T��(�ʊb
����>�Z����~��G?N�q���o�Ή�MK,���Ot$Ću��j��q?&볟��������r�`y��~��w���[y ,�G����dR�_�@��,�I�:�@8I �bq����s�Y�r�i��}������?!4/��%N�f�)k(\����?8� ��9�y晃|����r�2j�h9a�t�qןq�)4oގ"B�@��⹖-?+�
i70mlݒEM	a$��d�w���ݎ>��c���_/ᏜH�a|�+_9��/���KNwB%��"�5A x�������κ�?�j�h)a<��s����{|���Z��+5�>��w�5�	b#�⍬�t�^���H@H���t��O��s��i3&�����4��$����L^��%K����vۭ5f��0.���?����B���j��ƺ%+b0Z�p��'�e2._���}�s�Y_����Q���_��'�l�$�h�����-3�[JW]}�	7�t��=�V�9E�w$���R�U)Z�`[)ל�j)a\y���$W_}��4	㩧����=�n���;f)ŴYG�)�3QA����}��ٳ��|��ߟ�{k���Yok�!o��④���Θ={6������6��ʛ�c$�����s��丆u��w���~���������`%&���"�E�'�x�Zqݖ��z�#|�p�χ��(�ٸ�b��9�ݬ�a�
�,�ŋ�e��`%o�scJ��\��w��ElOO���'''�Q�eaX��b��R܈^t�A��CصU���|;��ΫV��@<��cq�i�5[FO�����9waÆ�o!=1O7���''X�Cs�8�9s���gvn��V�X�GBo��Römѩ@�K�.ݱeץ�cƌr��`��6E�Y��&n�vp9@<��N��ݴz��Zu��^{mF��zk�D���\�r����n�k4����n���v�A	�ʳ���Y8�r�I�1���3Zu���y���	CɾM��L|D���I�ܻ����fx��&�fs�&+a ����m���B�44�u<I�8u"RxN&�����e����(��0h+�u����M���{����I<ĘDb$��y��f�ey���,:F�Di+G�y��l&�ɇ��,�Z5ZnK&hnِI�~ɢ�� ]C������G�\t8�@��c$��pQS(�b���dA��fc��|f�@�1"[[�4�AFK&�RQyE1��5���
����300H��J̈́*�O �	W�8��H�����?1<����Ds�K���2+-�}�hp����f�ϙ8��3o}c}����\=�붌0���Z�!#�-8�4���A�@8q�v�����^.��.gC���9���r��	�ɐ�$�0 =��,˥B�P�c�%�#�$
�h#��l�ha�p�+��P)�d�-�n���E��b�,�q,�cK/p�;OVrVK��q ���4�<�!�`n!��rU�pŃh'1�To�s&9��$�J����i�ò��G�iG���pY��J%l�ǜ�䵵A0�6���@�=��N�)�O���;;��B��){Z�D��g����9xUIIĕ���ʥ���N�9'��9ژt���D,�)r�J@:�E]
1�F�o ���c�Kϟo��_��;�h�5�6�`D3�T��{"�p�iӧ�?��:�5%�ϻa=�S�d��-�-�1�'@�mSM$.rȾ�����|;��|��fϞ]?��w]s���9q��xԑ�w�GN���;�8ꨣ*,\^p[�nV�8X�/��ne�F��D2�ň�Mx��t�mw�׾��2�����p���W�"	H[s`���[r Z�c���ğjU�=t�O��m7�U�t3��4>�K?vʩ���k�������~�/���}h���{�;��v?&�4+���=������7�y��@���ض#�H�8o:�pL6'W2Z�i���&k�*qpHM�G��_͋��,:v��W�.~����¯��7��v=�����8�?�o��Ƅq�㤎�5�/)�9L�n`?�tJ�D�����f�6)ul@rj�i;�/��8��aۺp�O�-�e�Ϋo�麅�v���+���/���1������ʆa�`�$u4p'�d�Ԣ�-�N�g2�|	��d���c��W	.b�h��~3�h�X��������q��_[�^��/ް�N;�:��!-�Gn�V����c`4ńZr�͇��)�dd������;�v�u?y�G?vƒ���g}�/�4o���Oc�������;bƮ�5�p�U�!�}$���%`�W�a�7w�r�/��r��xξw�}��]��/��?劯~��Oo��дz��L(��BVV�M<�8Fw+���	#����s���=������Ww���;��e��Ѭ*\��u;I8���u����%�`����1��m�}�{�\r޹�]��.�={�eW���oY������1�b���%~�@�*�?0&��1}C��'?��3>�i��?�J�6
,>v�����u�ǎ�N(����ئ�@���ͦ�~=I9��������0�/�����s�����Cl��L���PTA|�u0�ZEbu-�7%a4ڙ|�!�F�W,�0ů0�~��#�f��a��'�p��Sn���w.\x����ͯ��l֚l�)��?���%�.�a[0�:�rW�S'{M>��5y��?9s��#�Ng�V�Z��o~�۷^x�E�IE��
s��խ��shp�֪�1�6Y1��x'��~�����A����.��9p�8�1��JW�Y��c�r4��&�X�=�9F���Oj��s����s���=�<󌫘����ȡ�������<�OB���9��0��D���G�͜9s���5�;����n9s������)V3��M��F�_$DӼc3r]�b�i����}���p]�*����n{<��7�Xr�Fͮ�̥E#^7�n��[9ZKʌ%
�y�<O��bq�����M�z�u��l�o���F�VϘ��dN��m��ZB9E�1Ls�V�PEl�g��9�m��.L,@�nR�'��ko�w�̖��d�$Y��N��Y�2�2��);_�1Fw�01���Z�㴮�ũ���e˖e�I��~�'�R6��Ea�:�C��δS�7��sX�R)�OW�ߣ��[������3�<=�Ѓ�����a��0�D$�E�b�?�R�Bm��F��ߴ�%
UK��8����������k��RƧ>��k_��SN���SNy��]���o������D�*���Ȓ��0&��3�o��V��R��^uC����oe���対��Q�}�����NZ�ti��;�8nqk`j"�)s.I<�5�MǞm+[=6��e�qI�]�,tH�Q������E�_�S�Rؘ*oZ��0Y�S�_�٥���?w���y�G�������s�����b��re�` Ҕ�S��M�M�16��L.� �@nj&���d��"a跿}d��~��Z;�BVG#����Bt�i��p�����?�~�d|���G��bT�������1g�Li�500 �o�m���Z��e�]�p�%�Ă}cS��x�)���'�J��A��f�1T�WZk"������\�믿
�DU���@.{���HED5�u�*�EIh�������ъ�C�}��-�@�R���䮩�b�������A��
�a{{A��_
,&�䁠�	~?����z�>2�E�d�7e��IŜ���*��ۻV�%%�@���(��fh`܊봮p
�$/��v�$�K�'���Hg$ҟ1�j�ƍ���˚��(�0�p���5�؍��0WenL$�\���	�8��c4�1�S��jPK��~;Q�uO8�1�J���h����8���8~����`&�k�U�u�!�>�ĸ)R��c�j���)x=���uK��Vr���I1`";���̶'Al�oܦ���ٔ�k�o$z�By�ιNKJ�LF�h�WM���uG�Ҟg�>��0l�YՊ+�-���O"<�~=��U�o��#�h�Z^�>�c��Sa���cL�X�dQļ�-9�X�x���-�Veܵ� l�^����L���X��Y��Wl�h���s�d�+Y�¤s�� �N;�v2I�Os��78����
è%�d2�f����i{{�@+�;a¸������ř�>��<�(�j2Yq�o)te�\Τ�����~��ex`�6a\|��Z�j���^{�<<[���':����UW]u��>���o_�`��M��	�#�Xj;Ԩ=��pR�@d󛬣ӦN�J���B8�?����p��_�c�׹�;N`>�T$?��{<��*�-�܃|{��C���#���?���i��0C	���8�t&�/7��,�>Dzz�!�7�8�+��leSn�H�:a��$��$:���P(��Ƅ	�Z��(�b�{'�K��
�o�N o8�Ht��cpp�mS��Nr:'�� �JUBMz^�D��&`C�rH�q�R�\.	xk�4@�X��k�x���r�f�Y�(�[�2I��V��'LȎ0:�<��@:)�R�,S�M@�^_�]�1i��Ġ�F��[�ӗFI&%�L�HI��tOE��e���D�1h��1�@�J������iH�#Al ]g$����0��O�t�ϲ�U�'��1,��@L�EO�\�%����	�sM����w7����,@ {ǟ�ST�BJ���}J��3?�,N�s������HH����wS9�����\�s�ąw�YoX���&�a����&?K����D���g����#���)ND?�*�)Su��b�'�3��L�;�ǡW�S����:H���xA�`�a}B��'L�m�N�u�������2i2� ��g��d6�c��	�f�!ʘ)�{ȟ�MaP�Uf��R�n���ɷl�XS�w.��_�f�đ"�Q8F�"z,e��'�I�Q(VM����G����uV��V�R|6Bз
���xD)��a��cC��M��Z���.�X�0�`���Pd?�C��a�:���EB�O�0�8�>����l~J*��j�Sh��3x�[)?��v�ƺ��N	�gx�"^�J�L�c�x`��0�+�O\��:,�׷�I�*Lm��̘�*��e&�����:>�`̵����Z1��e��aa`x�n��i�j���<0$��P��q�S�x�@��d���ab�ۓW�2��	�e�vT�Lc�p�g�͟*g̺�W�L�$�0a\�݋�����|�s)'���Z���d���~z������_�P�^ه�"k!4�����e�[��^`���:`�[5��&ˈ�}�&Fd�S����a��hC�D�k9�m��n�F�U��2�D��,�4��BoQ�^����C_���ڔ�|���O��''c�3V�Cx�s�]{-}����ț+�`����\8���+�h=����++���������|����Ь^�����+_U�}&5^��yU�_8�4�1a�8���y|�������rՊ���N�M}���'?��<�����[�CF�Ȼ�������p/M��5cƋ/�Y]�-E:��(���ul���,5$7cF[��[4���#�X�ݫ�Z�:��k>1����V�~Xd!Ϝ!8��&Q`T*7�s*�T'����a8�N[:AնxU�-vg�R���g	1�ޠ9'��y�rW�^K�Лc��k���J�8�2���yQ*��avEp[~���o��Lyh��2�N+��]��SO>��1���ʹ"/m�N:��N��u���o���z#������&<�|⫞�5��a6���i���cPkPF�[�0l;��e�2�Y���E����~߈�]���Ӱ��(2*�遨�S,v��I��������l�a�2���A4�e�6&[6�Ҵgm�1�0n��?�;�����:u�df���%N��<6��5����AZe�������wڐ�E5��c*�����Yfª8*6�{�:n"#e�3FD���15�f��K���Ղm
�TM}������B���H%Ū�;N��xm�>V�q<�Ib��f�v=2~z��~��j�H{��^s��7�ڊ�������]uH͇�{vY��ӴE^Y<Ł�=�Rۜ ��+�� �5n�7z�7F��l�1�]z�7?������O#�/N��q[��'��s3��&��1���t�)�GFF�����(ӂɏQǣ�l����:r���L;��^s��6yٖ�ڎ���sh��������>Y��Q��m�o��T(l�m�{��]�2�,�a�ෞ�e���J`K�cID7
׍!P뇬��\ެ�N����j��/��y�5p4��>�v=��΁0GE�c�v�1-�@����۳���(�e��ݨ�{�r�Ƌ<�۴׉;0��]��H!��M{6	,����
�A�ӑ����y�в!�R�y
����:'�`k�0e�qVN�6��z8���1���9�C�
a](d�Q�Lo�V*9��08p$3Q��4����<~�i��R���*Q���M�ԫ�O�;�����l+�E��0����5>-q�����.��h�.;�`��`e�ژ[�\�VU�{��S��R�����G$�v�ܝ2�IAy��R/Q���Y�y����e�yU�8�E�De��jmE�&F.\��ڱ���pb'O|�뼉v��7�9���Z��z��[��$�a	�p���K+�Ӯs����p�������P�_O��/�ܗ�A�]Z��E��TIt6�l��l��LhU������������p㭉������yÝ�M%6��TF����ub�H��z�H5w6Kܜx8�z������,����A}�=�LEU*�j��6�9M�"�?���akǕ.�&��}l(�APhR/�G�bA��iȿR�'�=��I�=���UQ�$�A⼍A�!��x�^�F�+ejgkg��D�gH&?�K�O��(*Ih��>?�_���PY�V��o�� N]lɬ��aȵ���R��<d��L�� ������FיS֘`�8>��e
m����2��^�~�}y�u�oh�,�01��L�Q*����ג��S?�bŘC��f�cJ�0���Iq�d�m�R�F��ވ�e���(�����"�%?m���]B�(G :�	�4��g�-O�R?�%B�� �hC�7��,�l҈=F���ұ@�G�
�#0a�g�̚󹙔�����	i�0�6"��X��ux��������ƈ�2F��U=1�R��O]v̧Y�P�;�?�A�d]b5مN&��{;��NN6Es+K�PVd�V��m�_��=�}�T	ҁ\+`�� b6�z����� .'��  T?+=�g�������r)
�a&eD�j��`q�C��D���qX��+�Y`�e�XD8F�O�"-��wl�~Z�6D�2�E��&/�̈́P���N�ya��!6f:�(��Ї�7̒�`H(*�f�XBw- �d�� L�ejc%���b��/%<^�E�����KT��M7vRi96�P����ׂ�����%�ʴ��R�t
�R�qP.�F�؇�7�y&e�GT4�� JF �G�����`����+��,X4~�]���l�͗0M��K�h�&�v��)�����x��L*��>X4C�
;)�^#r�<_���o?��h`�� AVȊZ�#VH����5h"����w"�G�χK�]�Akʒ�p�y,F|�T,f�>��1���+zP�D�C�d��"�L� ���L���X;,ZB_�"�!�m���3��I��2�tA��D�
0�V�b��9EԄA25GQ8sɄ�BJG�� ��e�?�)�J�]�����X"�J��|QF-��.�j���0D$�S>/�
>�7d!Գ(U�l,�0�J�r@��<bšDgRt3�����q�r�M�F�T����[�S��V��;�&%n���6���Ĉ���G��^4yc�Ԉ��6�$���(�6-�\H'�p��P�
�MWēMUb ����WFT$��m=m6>D_/䟞(%���D�Hq9C�|%>#э�rMj��P�91�y���#���{C�Ew
c��"�_���ޘ��|���3R8E�(�.�Cs:\_�|Yej��cXcG
3�5�Dk��^djq����;�R%��0�ݑ(�"!��9��P���'�D�C��W�/�J_��{$�(9���,�G$,�l&�	W?T�b�sX��
y�9e�B�
�iQB��}�ܲ��`��1��Q}O��8�|���(�0�c�F��(W��:5�Zdَbq��WT�v�T}�g��}@/*`G�՛Ĳ4ʊ��Uiu�;p��5C�e��D�	X�����	&��(9��f��p�^�H+�X�HqAc��J��4��v��H�[�8�1��>�d�����G�m�,�S�u'�>b�����BP�q}�R�5SDф�|V���x�.j�#6�M-�#q�Í��F��5�U�]�+�M�/L&(1g�������������X�bs.L)	����(�b7�[�2��B�ն�;��w�S$�Ѱ��~�h�T�,��<�Ta�_�
�{SX����8 n~����7#�,d(�4�h�4ŬS;
[�����xN3���"�E��j�ǉ�9�a��8Ƹn�(pvf��7�T�b���Q�Y�ld)U�PրUi�Y���bd�1��8���x��q�k(=A�%W�.N�9@鸇��6��6�H�~"1_�=\���&�и6a@y��3�\l��&��GyT%42��`�q0ڢ!�`]�b�ITi��xp�0O%�n��[X��Ӵ�G8m�1��q��NciKqb����	c\#VR���@�66��g�����O�� ea�D�(d��q�dL�K�&����/>���b�6s��J�T��UWe #��w�*�v�4d�4e%4N�F��L	���XU뺎��*:1�� g���i�h�9Hy��sfQ��$`�cS��aJ<@�a�邖���%bK�h�ڃ5��5��X�-�s�����#�g�Y�0aq7�{&0 I6N�8�bļ�,Y �f�E�B৞�z�Q��t�OJ�Mg�Ao`����Y��<�ê� ���������Ar��^��!�� ��'mJ����2q���sT�2�@��K����(�-��9�	,,�D��4k�:�<�2�4��I��< �: 8sr���T3�;�c����fnQ���i�[}�e����"B�j���w�b��mJ,V=;�&{�Z�Mִ�@F8�R=�aċ��J�.S�]y~�6f�i������W'7��)S�O��DQ���m�PDQ���xd;���xK��d��A?�d�����+N$J_�(Fù���P��fã;�!q!'��������H�O�Kވ��"T=�JL����
|_&p+�'+,�����aQY��?��3���+�e��,X���O4�ﻶ8�&:�h�$��W�'ɤ���9�M�ޫ�rh�e�c�H��H$�XIq�b#��0qYQo LS+ ߫0����+�H�Xs'^�����e�\Wi9��i���I�E���$M��	8�T�8���F��� �jHWg��Qۜ�C���"��:�ق�Ļ�(mz���ɅŐ%J9��L��e+/0�ϊ<b����	�X(s�1R�g���$FICX1���@�c��,�W���=}T(��*�F�
��,o��� �j�)�0��1�ɫiժ�|BJb� �������R���7�o��Z{� �IT���$�u!6I���Sy�^[��A4��K��1qx�:�9C/K��	ϟbQ�fh�LY�2_�.��:�N���(�#�f�N3����>�Hq�!Kt�(gieSG*C�ę���@,�b�����,�"�&�cK��F����UQe��㇅�Jj-���;�#�Y����W(�1A�9*ȸ)����;h(J�uR��X_�q����wS;�D�h$!oڀs*`�XW�5����l����O��sur&���Rm4�{��,�||��2hwQ��x>X�j��!�'�A��J�T*�y&�
�_�bT�c6�� J��1�'Fb�Xm�#*� /@�����4C^,�x9,V:�[%yRBA��X����	��Z�,k�a�5r�a����]1a���ڌ�tl'A<���iPܘ��}��t"Oղi0.(���q���!$y�E&�
s7q剗��P�]��\�N�_�����N��>d��C�X�*���� �o��&�Ԭ=���YN�<v�I"ǋ�:ZL.�j7j��m1�P��7S�6�S���r9��g&d���Krt�z�-`B>M��i����/1q�
��f��9֮s�Q�aa��FcP�L�����s<ǩ"&�&]�V�C�R3i��Aui�w��$��_�TYl�G�%L��c�e�N�)����}�,> �)��0��z!RO��56QbF�V@��i�1'OE֜ײ������s���ryuX��]_��ꄋ���^���*�;�l۲��>E=QAN[��XD �v����(�ǒ9��9��N	H�CQJ��<���F���	Ew	"�1aDl��R���Y�xc#�Zz�.�]L�Y����{2W�dR��fѐ�c������k�#�ֳh�W��Úc��G��D�&쨋��h=ǈt��j��)��Yc��'ކYa��~����L�U���@S��.3G���8iz%��o�	Wx+QM�O�9��Ma�s! }"�P���	#�,[��\
�T��"�Ֆ���32$Fo����x7S:��f"B#��b���u��>�F�:EA�0 ��u� )����(����U�_N�oX�QJ+��j=d��#��ۈ*�ߘ��U51��ŏ���2J�K�������ʬj��M�I�\�I���F .���zVEW��H]�H�F1��]��j�Ni��u�GM!�
b�/	T�U棸J,
ewF�x/Ԡg�pr�MQ�~���§��8u�W>�H=h(1I�B2��b�a�U�C!���0�8��L��= L=��5��&J�5��G	�N���t�ر������2���c
�K��]�K%)����^���rRH.S�bI��aE�"��Dj�L|�����Ig�ћ$M"V�6��� 55Ľ�Xob<B���3�1�B�u��g�5R�	_j��G#3���&!*xK��c�J4�h����$�@�{_��u���RJD�<�OLlDԌAR�K�B��j#"Smr�)4~.�HGx�i�@L�d�k�i����e����hXE�Òg�@#��"3�֐�`���¶N۰5��z�T>73�HF�s$�������J94����������a�a�cWU�� CgV�-�G�hK����6�c��9'��ǖ�M𼂫h�7�Ok�(C�.�M�Ex�r�)`��TF�4D!A���Ñ2UVL���%�BHEmC�)�J$vMPǰ���ݫج��vA`�á"- Ԃ�fɡV��u�-Pe>�B�x�n.�xf��@e�+(P�;��fJ`"B*��RJ���R�l�&z���@����:J�]�~}E4��E�w��|&U�-��s�Ɏ96D۬�$6��]�la�n��%2U��V��g�d��H��,Ca.BC��f�'p���@R��Vk5�]^ac�K�/�7��4C��" �%b�R1QD.��&���r=��|�8#�l��gR>[sE�Fl���:�9��G�ceu�C�� b-zH�*F���'��6	�3��6��uٮ���H>����QO����OB�tq�H@>��T|�]b�=��Q�[��K	�R���~C�Vt�0)3I�Y���ua+.c4�9��G��H/�Dt$�*��<�5	?�!bn���5��'�X�0�cC�������_]��U]JB��Pu*��'�~�ծ�C���C%*2���i�s�CQ�Ė��W of
KV-Q\-����g��p��@��P5�ee��بD#h`*c��K��Td�P"I<��b��\���馩ce(���U��YA��6�Y�9Y������r�� ��^�\�@�rI�c]Х�����t���|��m�i�	�75�GV<"�m��)R#3�K�xQw�;�-��������L�Hsg̢:9�3R�R�����ry�"��T;��p'^NW)���i�c�!{���w��uk������U��Ux�r�i�P7��c�)��ԙs9)�x��ixs��>�r�5��|�,���bţ0�Pn.[ ��VA
e�Y�dޥ��\�t�]\�N&+DЖM���NTJdY���Di�ζv���g�à��6�_ˇ���*���`�*�%�I�����ja�	cc�.I�x�b�Lg|?z�e�'�7P
������Y9{�fP��3�|ǟ��/�P��)���R�r�H��}팝��K3�6+ǚŮ���]������3�U�pTS�\*נx����R.��b�`�S:;��,xa8|��^@պ'Չ�s�Z�*��(�L�" �2b�gsm�;��5R���4���V���LA���v*R.D晋Ʈ4P*Q���JuO�7��2�<g�#�B*b��զ&��h=�����% `�o�#́�/jh.��57<G�y�L~o��3��3OڃY:@�W=A5�sYތH�Oc�&��A����e�Sɢ�5͞Ӭ��i��i4��#�u��D��5��L�u��a�`������6�������I�:�;�8T��y��������=��C]S
⓱b��������S-ɯ�T��ďA�j�ژ�Qq-�S̩�}�N>VS��w����+��)�E�P�Z�klvQҌ��U���T(�,>P�J�b�O@%v�hM�F��<
m�=����]��󎦽:��������Oh�L�����f*�]s�3��&N���g�C���V3[�@�4�4E�_�5����7���1�{��Ī�ۦS�u�����wҒ����;�F�z����^�ǖ,�߬�:+�(�]G@�Jo{�|�6�[�R���2�˫=��s���A����6��޵�n4�};Z��rzt�2ZSdn6c��F:�s�Ϗ>H��:�FE#Cw?��E^A��b�*9�/eM���;�=�@��	c>�2��$�2LV���cy�tC˱� wb�O5!Y�ev�V��%ϧ.6W�t,q���{�dyfO�z����TH���נR��U����B�$z�L��^��v���o{����_,"�0��2��3��ϡ}�a�Δ��Υ��w.�{�誟�KSXtt�N�s�NL5W�m>辍n[���0K�t�>�h�;�q��4�Ŝ飴]t�r���%T��m;��>w�,�ޟK'��?���h{�]�ɺ��}�mM�DԢ��K��C�jLS�X�o��u1�sR��xuCխ�ݩ��P����Þ����O=K�f�@eF
��TDَ<�q�+��_�N�6�˶���n�1+��n�~��(CCk_�?s<��D��@O/]EUՍ?L;���^T��*Ma֎�co�=EG��m������S[@�ٓ���K�����N#�+g|���O'��jƌ<�Ȁf���`G�&�Ǘ�x��.Ru���}���鵥���DN�j��D�ͫ�D�|��5�)�1���'&�%��8Nb��T�e6��gd�c�Cec'�J��.E�L�WV��j��rJU�>�߼�������މ���V��T���Ot�^�U+ג��A��p31�����=����)8��t��t����>���|���_)�wSG[��Ţg]A/��Y*t�(Up������Bއ����Rɤ���G��ȓ�ߖ�~�`���=w������~�`0my�ӦvRƝFC3�r]�T+�N:R�q��p;���g�a���.��t��С{̡�|��W6�7����>�gr;w��U@�6[=�H$Ш�P�D_Z^e���h����H<��M���T���c&c�-rT_��,>}#���K'���t���oK����CV�2)��E�jm�X"��&�,��;�?��~������_!�}Gr]��̻aV�	�urbjZ�n��g��wn5h�C���}|;�cv�~��g�}j�fg���:���O� /��"Ųf��X`���=g������&������W���<��{������˾y
=�2s�_<NO=��ܮn��Y9�E��{eo?��S%9{���K˗	G�u�)R��ηK��g_x���v&��L�
�$�}�e�R�*	��;Q�vC�j�nc�4GUhA����C<�JG�y�$�ꬿ1�Jƍ���Nk�B��O��=_��6Ņ�*��zY�ɰY����>�	H������}����NL�_�yz�Q�Ko���A��LA�TI�R��葕颊��H�m����u}�����L�;�$č�zm�z�dQ�Γ_���ZCKW������f�B\b��������VV�}�ܛh���л�K��>��g���C=���)}}��Nz�C�C},��R��M�*���YJg34X,��`�:��"+�[gp�	�(�E�P�W�!�C�FO��=�Di�����,�H�(���[_i�[@���]�3R���VO�
�%��03���̲1i�tɝ:�V+���W�>���nt����1�?�[j�兒�5Xe��k�f��YNէ뮿��z�I4�Z��2)F��*��7�G~��t�G����ffS-T�.L�[W&�Jp���8)�'�*�*�f3a9y���ӭ�Wҭ����oٖ.:k�y��韮�9��uLgQӖ�� �M݆*}EVZۉi� @�V�؄-I�:9<�+�XgE<�fn���W��Т[��ſj8B$k�u�*cH삂��m)���@"k,e������g!,��_<a*�'��)��&"nqKN��e%U1���z�CA�ewz:���􁃷�SNؙ~��+R�=9�٬@�C��U�y����֮RT��>�@��˯��5��5D{�-��c��S{�@��O�7{6E�L9�(Y)��&��,[E�j/�Cm�5[(��@Zߚ54���?��O=F=����N�V3Kx�W��mK��so�颧�(W���#=PD�ݿ{�RLxq�� /W���1��L$�C>����pB1�"��L����R�0��4
.j�b��0b�{A���oF�['�W"8�並�*�@$�t2L �����L�G�Iz�C��R���H����|�?[����˶��7<E�|��t�GХW�GS�fP=����Ot�ns�c����DԻf�,����=w1��'�0�X�L�MW��t������s��ޗ�^�mfmO;��AW^�$�i�R>}3�d�Q-����T��9�O���Y;����h�w��I䱂�ڒ?S�����hG�W��˄m�ѿ�F��mK��z˜����>Ms�sz�M�����WXL�ie����X� bf��0'AV�ҋ�fPcˌ���d$Y=*4���*a�t<%��a��.�k)�16s5�6ݏ�S����$)EGU��zN�i� ѫ��t2�~z
=����f��LTO�iy碷�n��l.�؆�eJ�w�@�����
�|�4�f�c[*��'���_��=�2��N�ryz�%t��K���^:�sD4�ġ��Ѳ���A��
���Y})��ζ.�f���f���c��N9r�cޮ��S�_K�_��D����,�"Χ�^r}����C����'�f�r��k��w>Jv���c�;OO� Zœ�����S�4"�ď�RcV����ƪ4�I&���^(d�ш�*���!�	����F�%E	�3�S����.��`
T�M��s�J6���`��ѓ���w/b{{;�U�6���x�T������28eZ7[Lrn���֣~���L������`����g��B��V�C�C����=�)���W�be�����P��K��U�εI���`���^���>��{�k�j�nz`�tσ��D��NQ�Q��]X5�K��k��ϟ��n7���*��<�X2 �e����^��K^�+���ɢ�g_�;R ��JRyQx�(��.����+�N2O�hbH��e������p�&����g�~A�L���� �����S�PQWVP���uH�j�/	�>@	Hf��w���Q�!h�Fqp�P��FTc�5t;�$!��i�WA
CPS����)TD�8+���`_ޜ���b�L��,6��J	'B�ӻ����_���i;�[G���HY�q2�C�mn�#P��$�XJO�#��k,G>����p�Ä���!��ܬ�d �{K��b�l��3V����4x(�b�O���aB��Gg�t����@��q�p��o�v/�k"�
�S���ME9�5/}_`.���B��À	�C�'9]"�,S����P�[ .*�,-m
���*�WbK()m���A�=�m�+b�s��B`{��Ҩ�㤔R͛�+�F�g?	3�����������
Ѻ��<�X�%��B(=���ʉba�l�j�l]��a����*.p�=c���Y�'&VR�-䚘�n�
,���_�V�RA�H}2�GUAccI Nc!��U��G�e��J@��7�AJ?M�O�@���T=T�A��T
EN|i!)�Qc��P7(.����Cĕ)�{2�Ȗ������n��Mq/��#�%a��s1���"���b��(�^�RU��������� ��!PB�-��,Sk�MJ��!�rb�5' ��p�T�J����Zj����G�A[���yҗ�?���QT�ut5�WY|�'�<��/�k;��0�y1@��U�S���wL��NDo9a[�п��yA�@��*a9�eE�/R��Q����X�6�t"g�)Ś���V��/�`��'R�l$ʲI�Y^ &D�!@8 Ѡ{uʲ�$ռX
Jy���l��5\�y���8�R@N��8�9(Ub��3�V����0��t�s�
��d�mR����8�XԘn�P��V��51E�Y�x�� ��͵���<�����T
]Ή��pe]��]pٔ�P�֕ �X<�K���<���(
�b���yUI�����C� 5��U���	`�+tba��	��v�R�+��,��eQ���	��h��I��@�����ErA�<�j��rA<ӑT��-&$p+�l�.��M: �D.��1� ���LmF�C���!��݉�`���	��@8�ͬޯ�s�r��t@2T��@O��a�5 �
O�*�T����e3қb�R~X1��@2oul��\>��t#I�,y�A��٬bV�PJ���׵�(��6{FG�8Y9ˣ�W�P��*�_���f҂R
�jC�h� ����8�N�ιT���IʋfI�;X�S`�Pz�E�{��L&(xUQ|%��*W� !@�\p� �w6!�)����s1,0�[&B�yl+�,����Tx��[$Y�!0���y}͛
L)����!g�n������,:@U�O�*}+�//�bsHǄ��e̛��k�G���*��<Wg:M�>�� R����gB˸!�X'q��4��%�mTS�@w|B�^�s]�H}Op|��v�ڶ��(�Tc=��=��1J��1���U#��+7^I�Dk���$`(]@C��A$�
�w4��mw��Ա��T\�Q�*$������釩��Ս�0�+T�.��U�V�-�l!̢]�؎��4Q! .^�s��O�-�5��x?��TH�*u�G���z�#s�&;�N����̳V�����]�C/>��'���ST�~K圲|ϰ�8F5u}��#p�}h��?C%t(w��D�c"��x���??I�������v�K���!uN��5P��/���?w!��n�i�������A�o���@���g~��e�����(�0XT��-�4��L&G�����IauP���l�y�!�A�'�v�9��y���
��{���B��N�QřT�'�レW������_,�c����\CJ&�L�Pl��#^�iوf�;�v�1�Y�R��k��9�)���Eǭ��AO,롔W!�S��<s�|�u���\L��wo:e���5m�A�ʞ�,��3Xl�T�n��b���s��l���e��0���Ru�������fNTa�H�/b��h�DA.27~�5t�od�X�����'}�bS�3"~�'��1�5�E��\���6D�n,09'@[&պ
� �D4��giv;��� �Ѽ�	�w�芹�O!��Q[.m�������󑥓yP#�9�\�)Lp]i���*���7|D)E�;�i�	������+�E��iR��Y�E
���H~2���x���# i*�ZET{����M{��Ւ������b���b��כ��� n���q!��q�c�YA.�/�k���^#�Q#ҡt�cBj��F���*K��|�����pC�Ft���kؔ�H꧅��}��iC�e�uO��@�fٌ�E�2��{6��rq���4���3a��|���AJB�p �ԅ�&f�_3���&I���9�p�C�ur"#V�Z�� rB���$B�H�M�	���TX������%׍'u�F=P�bCu0lG5�&�R�R�M�+����q��|�8Pu� f��bԓ����F!:D��y�9N�)����
U44�k���5���yD��bh��-�_��÷�z��Q���~ �lE�ե�)C&�H7��m 6���cH G��(�v��L���-~~P$��R�����n�@��sǺ�f$VNzv�=���4t���2Y�W ��#
!kZ�����bV��L�)1W�r�4BK����gJ��##����瘽{��=� _��-���T�3y$���`H?�x�j]�d�\Z���J<��T�*�L�_I���t.��1p�2��=ߴ.�y����etKJ���{�:�M�Yʁ��߈Ԏ	<ޤf&�� l�*���}�ڵ�7����F��]�d@6By��,�8#�k8�$0��,�\I�'�(p�pU�$����K�Z�|���Hm8E)J�d�Rg�@�#I@B<:���T�"!vd���ä��@�Ռ���
C����J ��b*M�:��T�@E��GWrz-d��򘉠�x�̭`���)I 5?���Q�IٮqA��[8�Ⰱw�y'-^t�,8F6�j�~��E����˧�$�9m]$o��p�.^�.���
���:f ��iB�C�It���ZU�P`�H�_��T𹧞x�.|�/��N�J��}dQxA+v�WgQ�1�\ fE� .��"�^��sK�H�ܼ��H&rTsa$U�	�b
��z��]Ya1���Ɛ1\�UED#���(�?��ZJ�C��tEUX>lt�d��M��\P³&Y�9o�����5��%�!<�._Nk�RcS���q�r͆	
�){���]��c7Q�g��Q����^~��[Ջ��\%��~�4.��F,7|��R!2��¢�� �4ܲe�؊,�e��9� �NA�����i�+�C�T�PA�j|(�lGC�����ء����]R0=f��w��(��দ����a��Ǥ�[�,��T�$�Wzı���֧�s(�h�ƕ{`�c�ch}e�S���/7���C÷�:�&i!jd#`%�I}��l"�憱�!l|����7��-uC��b�I)�O)g���M��i�?��u95�>r�x��-�v7gش���t�q�aȦ&!p)0N� 7 ��=G7߷f8�~�ah�/8�'�8���~U��P}\��bC��J`Ѫ�}t��h]
i��n�f6,�&|�F�HQ2�lwY�jU60�\uBI���.RM[�H��}�D̤R���e��ͷO^�̵f�1��IZ����{:�3Ho�с>(���@�MD�noXA��'=�M�8<GC+¢�e�&�,4�Q��U,�()����d�|H��@�tD�F&Y�h���EJƽ./)nR)P��zS:Gi���T���b���+�F�
$��G%"{�j5N�p�X�G�ԼF^/f�����hː,r�g$'�AZ�l���=4T_5�u'�l���9�b%�ћ,�cP��O��zC)��q��M�Xx-�H��b��*�I\+�8,5��~*��V�VR�]B�Y�YI4�~����'8ҏ�DY�.����DJ���N=���L��Xz$l]m*563�UJ���aqE��d��6�q�Z��78�*����5�&�����Ł�:�(D��'�o�������:����A(�X��$��֩���br;�5G��i�u�HS�DFb�V�+)�I!�ULE\|r�tbQ�j�XR�Η�R��A���]R����|n�\�kl�jQ� wx�MK��_���F�"��Hİ�qZ�L]K'V�U~���|�:���0��Oƨ�����olA��S�E�tm��X�%f2D�IM�XNw�X���0�D�$AB�����7)
&iAb͑٤�5�X�r�H�q�J�׎�EL#=.ɻj��O<��-BE�5�'�
bڊ�%��F����b��0�M��#H8���/z2�eS�8N乮5ּß3�T��M;���Z8ĉ&@�@b�(����Nn�7^b=ڿ�|�GҬ���$��\�x	Qp������Es&���Yqn�|�5"�r�?#J��@�,�z[��@�Z
*a(΀^1D|F{mEq�_ƺy!� Z�|����4�Q��x��{��ـ��3}M�\�ډ���xƖԝ�8@�eDB�]�E��<)&�>�&�$Wץt:K�(%#���$nr��f?�'M����:�ǆ�a�s���~�+�r��ZO&�����M����D4��������f�~mD�%lisyx>�k8I�ў�X1��F��9#)�/(�f#"�ՒI��A��-5��X��5���ؔ��:I��Γ�=*b8!۳��L����bSߔX�/��0󖕇|�~뇆����8(3W~*�qC�S������3����[h��o�nh�=)��?D_}�K�S��Bۡ2���+V�A�5���[��W.ن����UOc �3���W �4��j������ت�$��_mW���'($g�hY��y�9��o"t����R,�u5m���l��wI��ύ�(��I�l)t�����I�H��:�ee�����q��rP$y5���>��8C!�%�,�7ְ�8P��Ke�cO���/^F�G�Uy���"�,�f�T���}������]��Im!I�������G�%UC�Ԙ �� �y1~��o�k��{2kub&�����Z�i��ZV��q.}���yC��	tP�L��� ذ�.ʼ���~�a����ӨR.�:&�~U�8W��+#e��������c`�D�2�Q�X���^we���G��:���t>h6^"�����3im� �ӷ/��D~����R;Rj�1a�wHFv��M��CC�(P��q��d��j&�Y*JP-A��A2U�����Te"�{��l�[ �:R�q�LS��-rR����s(䲴��QP#_��
^�z/�S
4��ç^�fT�&C�
b�/�@��K锋lR�yS�  �Ђ
���󔚳-}���h�\�t�cD�+�ӓ0�}O�@��8ڼq�.�o(�d�am����>�)ʙ��³	�#P�}�Ȧ]�Y�:����ԙ�P S@�i��zdk����#���qX%�+�@R����X��)}D�TֽPp��ՙ}cC0$�� �a�^�veG*�!kCu���Q�>M���-1� bº�<٬
�#��Uw�$�\E 4\�m�.p����!�P�sF2S�l��<�"��Yǔ؋�Ĉ���r֘;����$5Da�tB%j��d��=�|���I-H��*�-�n�z[D�� �Y���C�ֆE&�Z�����5�Ni��@�!pB�ZC74�z'	ϛ�*��V�T\��>�S
3�UA���
��)���Y� �am:���E6�Do�q�8l ,�i�]��a��, �ZI-	K�X��Ѵ]�y��{�U?�5�c�*/�a��Î��c	9�ir�4���(#�<�J�R���YY&B�9+�U�k�G��7�j(�r�(џ�������6�"T��+��"E��G�H����%�2HE$�7�xk���6`"o�0�[#ͺ9���2y)��0t��ʴ�Z�x����](�	������e)�e�Hl�Ʈ '��,VA
��Ϙɦ��pr �N��&�j| IP|� �C����AҸ�HR�IԵ�@��㴊^�VH��H� 3pS�/�X��r��{rr$����h�R~/a��H����\L[~5T:�'�A�JAL�ؒ�&X]Et�W���`��A;ɿ1�x� �Κi`�jŊ���{�[�U��
;�*Wu��PMGRC+ �(�p�>�
"���lT�\L�- ���%�D��n�s���\'���s��ϩSU�T5��}��+v�s�^{�9�s��? 6P���{������j4e
�� Gd��zm��tݼn�t���[@�.i)q6�0R��ܥ���	�Mم#m"�@�:+^C�xl����2!�����ma̜����J�,`,GS"��5� �\l����u��! W�\B�0�e�}"�p$���1HR�E�a�vN������H��S�o�R�A�K���d��bcЛ!��������إ�d����5,e=٫m��z\�ְ^_%��5�l-\���We�#|����O��2añz�\�
�S��p���VD��J�b;���v�u1�F5�,���J>�wi�BS�f�X��!���u�^(�U��He!�q�\�\����b�¡�߹J�m�AD����H�n4����v�Fq]��~o���6F��P�����������gMT~��螰{=�v>H{i�����{䋍��)<��/�6�d.�OCTkl�0�����g��U��}��U�Zް׌l`e����'�"��ᨅ�v�x�-\�l����#+�	����Ae���ρ�!�(Ҧ�����p���H桫;�R�nӊv��d�<�����L���+���%�XT����%?��=J�=+�<�K���I�F'�k/+�v�U��9��6?��}�Zg�*��[Q`�La�XeA;`O/V���U�;*yttȩ�q�/]!��U�"���tG��/Z ��@&BW�3��|9���Q�B_�F�-��X�Ќid�������2,O�.�!w�K�A�X]bd�Kaf#�ʀR��!�B*цQ6��q��ܴ0 t��U�A�:A�� �fcQX4�����)pH6Q���Y���y�]��i��.Ϣ��f* �nL-�v�%�]��ZMVJ����T�����l�,.LmC�,�'wQI��FS��_�8c��^Vny�Y�RL�GDAe�i5�5�W����p�0ϲ�<)̂���`��et��� 4J�><�1,	�6��)Ѐ��+>0s,���B�Y�m:AQuq��w��yV�oҎ�»i��*�`�vE0��'�ob�@����+-����"��L����H:F�_�"��mjC��\�{[�	��s=j�LG�!�BZx�z��8IՅ����.���Պ�]T��Ŭ9�ՙ��υ�}&����j��)�s��	(��UXw ��yMթ���؁μ�,i��PP���16���Za��U���X��������+���M]����(�o�pK�z_8�Z(åp�8<2��ƁұN4'{�_��)��ܒ��z��͒.�B��#S-I}��al��|�ν�

�͊��/8_�H[��.��>�,qU,��k7�3�Z��k�l�؄2�`H[�B��,k��y��T5AE@_'���I��m����	5zi��Н�Y1��3#
���<��f�F�}�;��L�����8�ź
8��C�ݑ��pz�b'���Zp���3o���[���1*����<F����-\f�}/�@εF%�Mb#� uc��}X��ݷ
�.D`5!�������G�\~�:��8�q���P�h�k5�.t�[>4��Ѣ��otR�s�	P��깎� {1���s_�,1NRY�s�ե�8���u� 3��֪����.SF���zt=�%*"v��PP�{�Ư(��5qWݼs$a�,集
,�P!��K�ّlKo����4��Y�gӧ�Wg���K����T>�3~|R~�ޫ��0�Q��XN ��˂�Gi�-97ͱ[h�U���`ߏ�j�	DY]f0>�&�XPL���\�AI�� ��|�C�|�v�Y .T�{�����[��Z�w���pж������5p��l��✹��Zs�9,r��!g|�
��7v�T�q�[H<�׀%�Giuu��PL(�TG�vY1�tn�,׶ �5w6�-1��q��~���7�n�=A���]�ɰ�%�UQL��?��ی[��������D���wcY��E7e�n�Ge��TaƲ�쮪t����:C6��J5hf�N5��@�����ӻ��j#4�5LF�wzd�w��r�Li�̭���`"�{鉱��(\ř~6T?�` ���**�V?��ĥ:�X%k q:kU�;}ͼ�Z������HS����}ZGr��!Υh�u�l�$YҬ%� �l��F�DE"���
��L.��X���@�x`�af���<�>�h����`�ff?�����A6t�^U�$
,:�e���a&x9L���bh�
��/�Ԡ��c�2���:�Y�`A�9��/��$a��硆l#n�2*�r��瞑ZX Q��QW�Y>�<�`�A�nQ�UH=Gܥ#��Q3bx�:��I���*�D��պL�����D���P�N�-��6�j�g����b\.��ws��2]�x�C�p�D�����C�G��%��pp�v^�8�yO�7��
0�la�]���!��Z��0C�x�WG�P���D�I��>��a%0��Tpa6���j:�қ���<�s/C�3��x���J�|�g�>s�΁!�C��~���}"��� u�-�)f0��`��X�1V3EH^W���Şu���ݕa��IbB��w�^�EB8��P�6ѐ��;�W�D�z��$�A72�@4Ks�z�|my�����Jn���%�����!�4!���WZ8(��iny�^�D�ZD���Yw���u����JS�� !�U"cĬ+mm�.��R	�
J
gZd��-3r
e4�4
�g�<!q���,���0�%.��dlTDd4���P����������P3�)Q�������j��������/w�F��6��?��r���b�G�%��l����`K$�I��eW�����\��7������������!�|;�>�v_���|�&.���!AA̼�l�O���%z$ϥ;L�Zv��t�V	���KQg�,�(��T
�\̾�y���~#�'�Z.[��W}6m�6�sM˻ ]
;+�@��
�}��f�9�f�G�j��1&�A���
4>�:�>�tSm�^q�B7+u��^p�mw�o��>Te�eH_5u�,^���zo�B(�bb���;����mh$�)4-�܋g�}�F�T�$*.��ۡN�W��-���,��.��Y�*v�y�\��
9��ݻ8ğ���0-����i#̓d6d�YS��Q�Q��w�43T��<-�{V�x���"DY�����OGd�q�0`�42���������Q4����ް��~������ŉU�m� ��pWDJ�ߎ٪��\U� 5:&�����T�a&i�Ҙ
/��̶���z�E�����~b4��/�E�Wg�R)_�ٛ+���5�C�7�ό�شc
�c&C�����Ǚ�6�s�U�E���2�-���aT��k(GU����'��T��F�`�o|��ȿ�Ux$3\�9&J劓����>�pn�]�	ga�1D ���9��N,��	>�8��HW��*�}�,�|�`��W�m�O�Xl��3 �bע��}�f�r���+�0�@��͊,L����{r�K2�K ��c���i1";�i����-/C�N�ZB���-9�d]Qrj�2�9N�&�H��̊���=�ϵ�4W��X+�G���0%�ݨO�{�n�v��6��#�in��$��5(
�?r���쇻H���E���1T>���Ԙ,�����6�g]!��}t������|O���Υ,�!��xJ-@5�"�*ɮ�z�+���'�S0ږ�΁½$��՛.f�3���"{C��I�B�}�>�X��ϋ��`h�ܣ��E�
�/h0�р��QXÒ,��K_�2[�>h�7�Uq�D[���l4�:�Z���ܠ�!F(�B����=����7��n��;�F����zzSvZ����fw���M���0L�T���Ȫ�#K���j�3��f��v��ڝ��wYp�G

6��c	� ��7d����^WR��2�hN͡GHC�����E0,��ʼ�US��(������5F�סU��R�)�
�X���*e�(_N�b�0f4.�>���Tm�HIIe���Нi^��M��&[���ɟך��~�\��w�Ei-��i��k���Sb�,n�<���F�sT���w��-�$�f1��s��4 �tM�Rr��b$uW����*��|��iw-���.�Ϋ�
��&��:53'�`�p2u�%#�!������ה��P���ke`�Kj�2��n����a�C��,�%�J
p�!u�W��P�$tY[U �Hw>^�cÓ������0�B�M�o�>	.�1��ݾO��!`� �1L�P�0\ڨ��r��ah�AUl"�ϒj�v�u1ִ��`=G/Z��f�����0�0��K�Q#�Q�ѓ�C��@��}:�=b��	�Y��\f+�Wt:��0�PC4좑�P4�p�Tu����,��@p͚�ϑ���a��r�n�|j�Vj^�>�X]0��T�;	]��ik����;�:�p9�xB�qu��C�'�Da�պ�0FCw�裨�������	��x%6B��ev Z�뿎Żn�x	��>tn��y��X諺U�0��ynGq����ð�I1��;o�[���Z��j�Lե�s,�9}|�C�ð�F��*�{�s�Q�j���7X������׿���[s<[<�w�󝘒3T�?�Y6�Q��� W���݊~�t��#?����)���(\8��' �b�Z���s�v�DMͤ>��3�)�q�h�5�F]��p�5�B[dՄ�zwӒ�#c�ӊqt_KTv�O��v��ۀ� 6��\O����-c<�5aF�GVm
�[�c4b�E_��W��K�ߊ>P�G��=���W�0�5��nY���Pc�I�d�k�{�]s�w5��[���'?����"��������ǩ��0+��6Q�fk���5�a�qQ��%�&8��c!�o��@	N�1I'!/W��(lyc�Q�<K���^'=68H�qA�B~���0���ep�
d�Պ%ȝ!�X>��i	�Iu	��2����G����MEgD�g�A%�L���#�b('�,?�C�x\oԔ[�%o�LfM/��g�NL$�W� o����F�F-W��A����z�P�����:�CW8��'�l��ԁ��p[��ŧ��1��,7�f>W���J��J0a��i�c0_��p�9\3h`1w2��/��X��Ɛ��!�e������G�����͉�E���\�z<��;��� Y�2L����<`3��+��+]ݴ��n�s1~Vj&���BSs�D:���� ��!��"��D{Ք���+y�ۑ�H��X�4PF��A^X'��OF�$�(���9��rNj�ɲF��^���a�,L��>sJ�\%>�6���H�Pj+~�J��-\J8��s�*�d*����!{lt���$T��d,�K�����v&�n��R�Z."�Mt?X����\^&���5bEV��H��G�T/#�ˣ�O��c<��h�m�-��lsЩ,�
|
��N}��qҞ�\V��F-�v������F�%,C)�j+���tz_�s����E��=��R�j�0S�si��l�[4��eyc?���Zv�%y����l�0i�\�Y%����p�ى��^��uW&���3����m4�Se4d��j��r��\�ء����׮���������XHá��W��9��r�3b�u�7~@ꈀ��U�s�p����i��3�z-���\�F%����Hܢ�(�W�ԹID���$0ʊ�0�Ct�*6?c6�V?jq�����䮖�ԁ��y�P{�QrG儮f5O�jy�8?����劣�cC|ٟ�/��V��u��:�YK�4���p�d������B��b�����zf���>��3�׺������h�lҠ^��f�S���*Vh��C]dj���!,,�Ccj��h�kDXL�$�z��=�Z�J[	w�K��P���]��13�p�uX8�X,���+wlP��`�Z���X�xbT�:b���a�bLD �a��'�@ֶ�z��6Xոb|wĀ'�wsfN�K�b����Q�k?�#�[��[��.�$��F�k���Z��`�#�� �O��fU�b�V����O��d��M8���H��X٢���f�J�#N��B�ZeZ���μ�"T�ieVL���Q�0��=�����D��AY%cS��A��P�S�qR��5�ﰿ�ܪ�iH�=�B��3��W��/*�͋�ُ{���oV��[�0�q'6nݩU�D�ٲu;��E�sF�Q��Ë��Cp��3l�n����a�����X�N��R��q�]D�]¶3��h�u5<��޽���_�+x���e�y�h9^f[b��p�w���}����s�05C(��QmlG_��bs�Y��Z35�����>Pv"c�����������`����'5�5k���{�`��p�����?���6�U�%.�d��G�.QwX��*��X,����{�w����;о�غ�Q�u�` ڦ֘B��]|�Y$b�(~W	}ߌS�$�50��*K�h��٬e��Cr�����2�ۮ�]����ڌj��ޔ܁ͧ��FA��p�9���5�Hs��o��G����5��3�}݀Ab-�A�2����$���G�	Z+���$#-3��:VP�1��e����p��ؼ�j�ɹ��[?�]7|��kO�G��AqMOd�dh57b4*�I2J���>����<Įͳ�=�sӗ����T,C;�Y��J��pB��R�2Nr��w��'9*��u;�VU��,�b����[����_��?v1���/��s����7݂g=���W��٭h���Q�"m3�?{��>�q�>�t��s������K.C�9����7��g0���	�ic�Қ�5E��2>��A�&j��_��C{P���/an�"��~��ֿ(d�7?��8��]hGm��]���|�tӍx��~oz�_cq� j�Z�6��uo§>�y�&��A��K�?7\w5��18���\`���5��?�J}Sr|՚-9b3@1Av�`�� �W1"7l���� ��!->|׷p�Eg���y��/�Қִ:�t��E�X.��|����g?oy�[�`�E(^����شq3Z�SZ�ڜe��H=��/�?f�؉�����'cnF��Զ# ����*|��r]'2V�DO�k���o�͠ڌ�_X@�x'���g]�{��y0���w���e�k
��n���]���/�Kq������=�T��]BF�(ǵ�݋G���q�/�<���{ދl����3P��&�����2�t�B�qJc��`�D-�`���H�:6NGX�� �q��.�K���g>K������s�t�mk�c�y��/~��睳K���DTd�%w�w�Kv����ڨ0'��?�����w�̳��\�T�2^8s�8Y{�sU��`����LqcZ���b� ُ��{p��b3�G苇��g�� ���û���Ӵ%!��}"�u�%���M
�Y"m'�V�bW�$B� ��oԞbc�� �s����P�R"m{��;w�x�ەl�k����S���%�r�
�9R]"!�r4���B6w�zأ���R�h�����g?_��y����(GG[<����#��h��Zo�,��7ߌ��/ğ��r�v`������.�o�q0���t�����(���O�g9����z����V{	ƂR8LgZ�J��$b~�0zK��P�g��x��]�L�,݃�-m���5���bt�\������'�u�����u�1.����܅�/����w-�E��"]v)�Ze��{�ޡ6G/_@%l�ݚFczڪ�
�q0��p�j���ˑ��T�kR[(敫�����()z�ƬW�<q��m$�k�����eg�Ш��s�]���06��!�i�u��WkX��Y.���L��&��A4�����P������J�(B�6i[$V�	1E8�t�be��)�q��`�E���#�*c�cܒ�5�$�CZhWW�;�f��ލ����E�,uPW$�PqA���/�u�zl<m¦�(DX���%��7��s7����/x�s18�u"7�e�aϡ�\o�μ�B�$�+y�0D��-��}# >ec��?J\9��g�UD�'Y�Ѱ��[eV�(����]���n?�n�zK["?����^�R4ڄ���h��7�WA�A������mÇ�}�d]<���m��#��;�ȽL#I����\õ�f��1�qq�b�e�Ȫ'đq�S��e#
-'�&J�a˔aHvj��g:[����}�k_����0]5\�/|�x��_����y�FYO���r�x�uZַ{�yj�Fu�N�眿��G�i���_Q��T_��7�8W�����g���v�]=��>�1�3
�Z8���:��� @俉��N~��eiQ^����p|�<��/~/{�+133��7!�E����q;�6o¥��_��c登��Ba'N;k#��m��v��>�ױ��a|�S�ö��������e(d�J+�I��G�����`gxnu#�	5�Ɏ�e���v��ߋ��r4E��[/����ϨF)~��/Ŗٍ����1,�J���n�NO�׾�5ر�\����]���ۍ١�nD�~fozǻ�ܼw��JK�Ȼ�� ��Ѫ�(`�A/�k���S��GqD�y9&k��"�j�H�4���+�'#L�7`�����;���/���z�4ds��֔�]�y�]������w�@��x�k_���J\s�wp���ik�p�G��FP��W�Vi.��_F�ލC��8�ZX�%p��0�v{�5�������\�uō���1فn�������ô���Qco�/�S����'��ϿQ]w�q'.<{7�K�8�� z����`��ͨ�ut�4��׿	O��_��7ށ3�:��y�D��0}�#EK��Ae��ulk�9x�
�D�j�����<�1t�X�I�d\�h��H�6@��j��im
�� ������c�;����o��ضm�x5�Om�:��--���o{3�x�p�m7�='�h��7s@�t�{��:bx��<	�偅:w]k@� 'S�ud�+?��p��eK`t�߭�1Ҹ��a_Q/&C7_AI���`��D��k�����x�{��v��~���Yt�0�f��3ӱ����Y�{!n�I\ӊh��s�c��qסEl:�t����	P�q��%�fS6���qJc��H:�Ө����,����f0�]�<Ksg��o|O;7�3�M�v�=�ᰂf��5���-"B$.�]`j�N��&�/��K�}K=��y�r�M�v���cv�,���xg����5�c��5����\]j����w{#eW&U����&"1,j lv�y�
9fq���;��$^���?y�><�<l&���{R&�O~�����3p��O��܅�hl�s-q���s=�l٩�}ڋ�	z\���Z��4F9ֲ˖�/�-���,�k�Ĩl6�O�Z^�����*GKv���3 ���WP,����@ܞ��{2�a"����1�s0
U+hLoD� ��c|Э�9�S��uO�3������7p������3���r�lFD�򤯋��"dX��޲i��,�gsl>�ǔc���3v*��2 ��X�{ϋ�*
�6�y�<߄F}�V�Ȉ��+\�^�XԒ�+%��/��������ʗ}�(?o�]����0��ϗ=k�3����_�&����6�1d�;2�sH���/���*Xw�~o���=�����(ĳ47���DUm�D���"�۷Ga��6�R6��&H�@N�K���+b����#l��F0�˄�V�T��KCT�R萄�2�U��A�I�	p�zc��5A-٧�Ȗ�$�F�7��n_d�:��~��ZQa�t�K4�������>��(�jJ�C�"����/�ǣ�0bT: �щ�\���ص+��D���*��ـ��H���I�����7��P�C����C�za)[�g]`�r2�d60E2IZj(��J� M�תW:���"�-��"5Ɔ����x��/�Q:�S�a�G5R8�@��=T�M�1%�y6BK��c�F�#�r�Qd]�,C>��>Eg��{�������6�/�}�����/���G��Ncl�4/�**�S����ˏ��WǄ7b�µBy�	@�b��exGUyXe$�L���=Z��]���I�Mrg,.Á�M�،�j����>��.
C�ue��|��#�+]��/�4x��j\��u4�R<;;�o�TQ�Q�D�<*Z󡛉��T�+���Mm�X		Gz�Xo�E�J��.��A4k#�q�5�֌l�)�S��ƍ;Ā��� ��FT�<�ZA���9����)[i$���/D����&5rZ�w���]FH��MA*�̣��Z���r�X��?F-��lT��zA�ץ��/�m��a,�P�_�M�D&m�hRt��V�����J�ԇ�X_�Z�X���b�|bG��x��P�Ȇr��9��W�`�T�f�`�Ar�C�؆UӟS��)*������u
`_�YZɽ��ĕO���y�]����k��M�[�Z�i��}����l�09�Z=2$�9wؖuQY}�Y�c閁���$\��f��5��O�d�G���Z�v�7�'�v
�?&�X��A*$�_�y�AODbńp������O��Kx��_߱(�p�Q���(�INdc�yi�W��rqn�E-o��D�[�LP1Ru�Yjb.�t������h�4yds��q��ɳ��e���Q��_w��tu���������e�P��5]�7��H��}��nwZ6�A;��Lz)���פ1��8��l�-7�X����UQ�Ia |�%#��%��[W�����w�H�g�`<�q�Rڬ�R:M���ڥ0U��3���v�$�i��d	?w�&�ɯ���'��h;�R���1��͡��.��9�q(����兯����(0q�x�=r(�99Y��T��UqS�*C4�yZ�-ٳE����!R[��[ɺ����}���B��[�Tɠ0H;x�/�,^�a��)Ɲb�.����Rɳ��A)�(�(C�Q�VQ8�l^����pUk.�X�?���\��1�s n���&�ŗK���h�t�f�,D�<��Ύ�J�a�:���@��N!J0�D-)�6�f3E�S�c�&�&���Xψ���������í�G��ޗRO��yZ����EV
ő¡~N8QT8\,��OP���8(I�u.�ٝ��3���P��CA�-1[�㮽�`��I�N4�Q(dÑ�%y�G��h]�@,���᠇��ѣG�e��*�M�L�b^�h�t`�C��nCv�?p�_J8]�I��t3���[������(nc0�x�K��)W�=��Z�'�����:�R��>�w\�s�>�3-�� ���t���Ck�9��[ŧ�������.<ː�s{��+�5�������� �p���D ��j,
�+RGD��5r�O$Z�P�d,��TwǎJ�kj?w<���f�zL�<�w־�Ȁ���نc�{����9d��0�o�:���hk;��:��b#M�30X����VÊ�V�Xa���jk��П@���1+36�����%����-�Xh����;�/�e��j<��y*����V������?O��<q��cœ��P�{����=yc��f|��+��>�7��qC�,�s��H�i<��+����~���ص�¯�ʯ�[�:���:���'xȣ��o���n>�#�UG�%qp�R��e
c+K����Dt���Rz1ˇ�'z�/�Y�Jǡ����!F�mPJl�J�`k�����}����'��]g?Y��D���*�E1�?�����{j�i12E�U�8q��5���,��*�w/�Z�`V���3��*�ܳZ2eZ��D
��]���V6�S̠��`wP���	m����n���,�XJ��p�Vh��(����Đ.;���O:9�bY�O��E�#N�"#5�*t�����^���)��F��"�F�C�5�YNG.�T� �P������J�(,�c�M�h�,�6�l~c�3ч�">��(I��,O2��������'��ۂ�X��o������0l�m����>�)�+[��8<�(Z���D�b?Zn~Z
�k�5��Ȯ+���G�o&��z"͙��h�b����C�s�u�Fb\�
����a�3��^�
���U�ᘞ��+˘��h���G"�5��f;�h��"��s6��\r�$@�h
��	ϣ����A#Y�^QE^o����Bc+�7
����|lj?7P������rI��J��1*;`dń���+\6־8\�y�[G��X��,�l�Ao��O!���`>�����6o�푙�Iv҈gG��Q�1��i�dRb(��AilҖK��D�9��P�b����gU��A��F2Pn����#6��6G�B�8� Oא�;��zD@�%=s����I�D,�sLM70/�e�X�$�"+Q����Y=�0�a-?�+�0��ī��q^Tk
�dN`krĈ�=����r������13<'C�f$��10��^K�w^ V
���=nΘ)F���.f[[1�9�ƝmY��y�|řh��ܠ�	���{8e��^X��dt՚�x�J��h�.Fk*��j
ݩ"@���x�6�T#��Ē�n���.
c"U��r�.A@�������@c2�#@#�/i<�F�yU��pc��-��Cr�1
k������\�%�v���&�=��#�h]�jx^s1�I/UK"������N��W��c.��e@�9 5X'��2P//��ɀXbЮ֓=I->��AqQE�'��իG�⣂̧�2h����&����r��즙Y1X���(j	�"(��l�dCl�{ZG"�K�	H~+�H�ʦB��
Y�D��������r<��eh��6:8(�l��G���|OE4G*Z�뢥�X�B�#l ��h�	R��H�~i�dnR��ж��V�3�%�s
�h5��SLe��ĖA�u���S������A��?1w�e;����QrBC�U��P�ͽ>�M��t^��	XD��\jm�0�C���O�ǣq�mP)�l���"e�������/�,l�[@�w��[��/NS�4 	�>
۸u���Ƭ�:i�Ա����%��IҤU[�z8g�n짶Hz�Rk8,�̉�PC-�Q$�<�����F#Nb?��U�X�{���b�ʭ���"�Qè��+a!L3�>�шvz���4Y�$0�&�2�Yi�JA8�`L�Q^��`Иn4���c��˼b�Ǣ�xlя��v:4�������-[eJ��p��()�?�aV�G9��8v;��	�L�ٕIĞ^�����t|ظ6n�����&�3#~��{x �;{������b;��g<N̪ȃm9���t&R��&M��/ޥj�,��f�^�|g��.A��NG��^�W��"��QPs|�EC�Ӛ~��q0Wk�QUW�8�G��}Ypf+C��(�]�F�-gwU<�@Y���⎒��L�	<���(2�Qs��=�%hb��#t�J�͗�raA4r�UU�WmY*���2Cz$�`��N�}��jr� �p.��Z�X�����8�b�{�����"-���$�h��!��vY���g�� \��?��!�N�[��J��� �L=�Bŀ:p��Y��?�!N:��qAA���E^����YK;����h�m6�_{Z1�^��x �ZZ��6W�2n�bw$�(�X��RO��b�k�"U�Ĵ�@���2��j�mlajX�,(��|��.\��de���%�V�P�3���9-ǤQ���%�F]V�#s��+��$��0S�D��Ȇ����,Z�`h�%-i�V�e��nte��D��-��]&�LŒ�ԵK�=��@]�x�A\���fԛ��W��gd�]���_��p�E�;e��C䨠��` �;�VE\�,��~����@��ކ�:��@�SC������	Y���p��h�� %�!`�
�)E�i�x��³(�,F�h4@�M��G��b�*�R�T���a�̆y��)%	�k�.����}+SQT��)�I�+��"r�����aE(� �b�����Y���xW5�™,�-�}�E�GM������yn��p,�b`���2uG���W��r�����8~�B#��4���ҵ�g+�" ���S�x��A�!�Hu٣IA�h�*6EC��"Ҙ�H[	y�e��scW�cQ�����+�ȃb�?��NTXp��b�G7U�4�IHEJ㙂�x�ުB�����!zWd��"^����(�m퓖ss�V��v�5h��p�H�s<�X�P�8�VܒO.�R扆��}��v�s�X�	wR���,�#^���S-��E�D�]�㸳G�Q�jq99��yD/D�!�4*.���q	߉�J���>H�5��w�r��5��hFa�I,��,6����Q8�\���q�VBd��zRdU�x�$o+p��Oȭ6�xc��:L�h�Ck"�$�S���Ƹ�H;1�SӚ�]�,�f��)dؽW3�|e܁@e�\�(5Tb1[U��bYeq��xz�Z�X�`��!�������$��8�1x$0��դ�Bn�(pVK�\�x��ʻ.�'A��6�=��1���A���Z��x���Z u�:��w�`��f0i�p��5 �K0\�^�����9P}�P��-�;$�6��*v��OML$Z=�~W�c��g�f/aK!G![�@'���{-�	�P�6U��rn��e�B_�q��	j���y���P�3����(B���#1�#CS�C��e�X#�h�t���o\��>J9Z1Ĝ|@*�6�ۊ���-֥�����Eq}�u᫟�\;o#�~g���/��̣-F%#�*8bwt��҇?n�X]fkD�Ϝע�:X�9=����]�>T�9#�N��'�e6�����E�u)�U&��8Tۤ��^-p�-�a��Of��A���"�zMÓ���u��Q�4�џ��M[d�&��C��w��ϽL<��z�i�6��Gj^���1ƪ������%�F�g_��~!ww�Es�K�z'����-���i�]Pm�П����p�Tf�k0;��v��X���,1��-��>KZ���U�Yո`ʅ�X��銊�dK^���5[H[&&��>���_Ʌ���(�R:��}��m�g�]��x�����/GO�d��d�����~
ؾ��6�'��K_{�֩,f^�8���dԣ�j���[O�U/�/^�2�6�@D29�?x&�?�g?�J۩�2��^�y�Lm�Q����_�_��'��h�7 �4q˾%��Wc����jaO�
T�G��5l\�����$��8�A!gK3��M3�X��7����G\����Qk��n�����n�\�+)Vy��5�ח<�I�͙a϶
j��~��E3U#��̆vY�KC�h����2N
�KK���}䪲#1�2����U�`{b=w��k+�B��[� ���Ɠ�������2�F��%i���u�#IG�G���B{%7�S�SF���B%yr�ꮲl@ٖs4*U+$�5e�f����T}��j��e�㗭Ze\a�Q�߿ҋ��%�EVVÛ��f`!���ES��H��9Y�,;���^����=���.������o�#���^��X��_)����7Y��2u�NhT�L�z�/D�����Ci�<3�GPZ�����ל��u���MvT�n�����ǆ�ѝ�Ul�l�dM;�f:�sW�r���5 g���Z6.�U�f�#K��]��xմz�aC����Ov ��x�2f��X�i�/�հ鍜�}a�e�{�uZU^�Ҽ!ih�8��J�G����c��	�����۞�o��o�uzX�R���Fk��+n(0�pƑih{�=HU�+��`<��f�'�2��D��7�B��T�pe�h��,�dWOq�C[��zR�86��j3���� ϗ.zY����.>B4�qBϑGG��*6F��-X�6��\���3B�[Ȉ��s��pe+���ɱ_}G�T|qn)%��I�����-������Ɖ
�FQ�wN����윂�D���V�[�����١s�=_�ڞۄ�s�;�q'(:#V���?V�1֮[-Wb����2ʨZ���{��S�6%��O���y��-7��+��WV��<�Iן�5�IL���;78�����z��qn�iP��լ��<w6�� 'c-�k�v_OC3��3K#>aS���
˝T5���G��u^��aBV _�� ���|p�dJ�C��]c�T0�^�ޙ}s2�K�Ń��3�%�h[�}U�c#!M��B��%���᛺���6��u+�(�	'~V�U��:�*7���=6��;�jh�G��;\�N9�8�}���7��0���bh�Q���|��sN�K��h�u�����l%YTKX�HT���(mP�:��+��݊@�D,a�Yq��F�y�(5�9������w�E�(Z��X��aeO��S�XAUo��uP�;�2��Lk跢���-v�l��e��&4���U%�?Y����Di���r�Qq�,+��,D��!���(�4�oB�r��_�_N�Z~?�/�)U7�I8� ͦ������̿-�<�k�"�]�ܮrH�YK�c�M�����(�)���e�Ga�Y�G�]��I�`��W� ��}�}��4�c��љ�<�w%5�Cd��4�����u���5�m�w��ǳ�����}v�z;�[ Ѭ���q�A������w�,L7�ǐk-�Ά��X��_#��l�(�� ��2���Ώ������P+�+)F}DVMA�Z?����ֻ��*4��i�NT�-�����0���,/���|��~��ZB�G�ח��$'uKqƃL�I�-�rN��1��(��(1�n�[y�z*YD,��r��s~W��Qva�"��h�M�ǲ�w{,�>���Q&����O^��m`��ziM༇�S�*'WY��_23Fc�Mkڊo��U`F��ベ���a2V1Ũ�E;�wؔ��Ga��^�v�Fd�&IZÜO�<`�Yl�A�>&[���� �7����Jo�w��+>�[�N �w�&�<L��������`�s-��U��"i~��!����A.G��,!]Y��΋�}��w11Q�V,�.�(\s".�MD�-=���m��d��jv�{(�й��]t��}'&j��-1��Pv���sx��������!O�
:d#U���b^��ui2�]������%,����2L{U��b���N�aZI�f��o:�_N�������c��ba)JQ�aMI���LU��L6��}�6pE�>����T�0ꃳ*e�����KP��;�X�T�βD�<*a�4�=�������>&����W.�^�%[��ܡ�X�#�*b�,��M���Qf��>��Z�jb���F�{U��Rg��+��=:r�d̪��i�v���}�C���
��+Ǒq� [���̝�'
����U���51���`��2.)�[%���Z�2Y�`1+��P��x k7iCd���o��zݎvw3�Ċv&�<܏G��I�;-�W<�������pYH���1Zǆ+6�0��j�JcF����:D'�jMk+r�īh�^��(o��>ܰ%��z�ݥv������Z�����Im�ͱ�
.mj^����la��\���̚��H���Jh�~���
ƭ�c���G)�f3�1��%pY ��u%�WLElMd2���Z�]����N.�/�5�c�����B�b�l��zl�[��!q�f��'�Y����c��E5d�����HG�?ʞa����i��q?j�]E[x^���X_�f�z�5��|�++����ވ�Y���':�6F�6�[E��EI�(tP[��U�D�S�:�y��n1ºz��e�~��p��K+�L���fD?�J���,�8�N�;;�Z��5|
VY��&�J<�td�
dD���ŝ8��]폰�{���9>+�u��AY�V�W�� Ř���}z~����.0'%�sS5Z��Gꪎ�q��C-2He���E+Vo0ޥ�$�U1�3Pau��XSd+&���4�R��ͬ�5tF�.�b�Vv�6	��T�KSm�]��z\�'��h���h
�E���r�[\��v�-6�&������Mc>֠�Q��EaU�
o���g؊}&�}�7��M(��GG�E���{ޕ�-��mP����y��cj'EiN������a��I3$���@1��tǛ��D��(��'2�$����d�5��U��E�^֘fV��F(N�h0�`Ҩ?R�B��,�Б�Ԙ9ʴ���i��H�LB�S�90ΨA)l6g>�vߎUl�����(�x@D����x�q��H��^}�@��|h;�g��(�[-�T�`XYs��D�xP��U�6�ar���!�O<��� w�"�r4vY���uВ3�a��ݪ��X�����;�&�|�f�1�F�q�s�?�fg��.Y,O��X�^^�X-W��o!�~��J�ɝj�������"�(��v��������]���6��*e���H��]�j��)G
���h���:�*��l��#�0NZ�)n����qF}�"��^����C�*�o5��ׄ@xOfbh@,�O�4ǘm-p%y6Af��k����4L~c��d��Ǉ�K�s�����e]�0��m�L�c�*��c��ǸgF�r&��~��F%6W���^g��k���C��/G��/j�k�5���f�M��ڮ6�Ѱ�Q��B����jL�+rx��
i�Mi���Q�.�gv��|������k0����������Ñ�� s���Y�8@-D��i�X��*J<���:BWk�,k��S��f��G�w0]I13a�]�����Y��k����i[q޹�cv�F\�5���7@�kϾλ���۱Y�%�-Z�1-�G���Pm������hh�r��r��������bBN��x��L����Iy%��Yۨ�	�j��qе�Du�S0�D1ĭ�� RN�I2��3���(��.w�Ot�H%��Ii	�6M��W�;������x�_~����ٴ˱z�^��$���V|������֕"YS���	;/}8n;��-;��Qo�����8��4A�q�iC�D�f%,r�I|j��ʚ�0\�D�7J��v��s�@�F�4��¥;���M8`Ho4*�����KbC]�1�[-5�r1�'
UƑH[�p!�X�V��\s����ѻ��q՛��z�c�
䣞���Y?�0=;��z�x����o����}���O�7~�٧�;8�8m*�-�0�b�����oEy�c�T��Dl����}Ѯ#ͯ����.()���_~��#���O�R����@�*b-%?��Ǎoz�|K`7��JW���Ko�����0�˞�r,UN�(n:��,76�a�y �A(F�ᥡxm�%$�Z����8��}�U��]��k?��wnr���թ��:��=d`�������?�?�����Y��F�L,�50Ԟ��:��&a!������]/8\��ڒb��a|卯uu �6;�|n�1�����bg��KQ�r��-2�H�bB1��kk��,��+������`�\����L�A#Ws�+���D����ȣ~�"saU'��v��tw��O��M�۵ �#���,�1�%�R�0�Z�T0מF֛�L��x��G���6b\=� �c_�_f����8d�����W��w��k��U���/�����Tis�ץ+�TE���@0��s�ծNe왠$���&�Ɓ�:W�}�ӱ{Ǵ�0^D,,.��`��  �:�����u�=ޅ����	��,.��,?|N4����:K'�@!������p��	`dq1���dQt��+�VbɤV�"di��S�aK�ŗ?��x؏?��P!&Vl�),�D�q���B �@ql%��ۿ�CK	���7��]��,|/]W
�}0ֆjE)��������T�Dh5�sS���X�$Y��j�1e�]mn���-.��"���K���˰�T�⚆À� �z�D�S�������+�6���d��,ʩB �F���gl�o������ܪE���Q��~�z-���(&>���!	[M�6y����|�3��~�|�s��O�|/GufZ\�B��x��d"��`y����3���R(�>;�"��W,]$.8��LOOc~~KKK�29<6�Ɏ����D+�Sf;�V��/N s���U��"@�{�^9ƕ��*!�}���1ը���V���w��� 65]<�I5lV�bJ@���G�����Ǩ�V:Ǐ~�ݯ�E>�=�hO��ngQ+��j� u��V����	-�c�!����E*\Wq&4�Yg��Zd0�(���f�]���녣�U����r�\�;vh�Dwq���H�$n,�6���w�]�y�'#ɓc^��lLo����Gr�d�{�5x�c?������Kt��0(�������2~����J��Z͚�W�B1b����ݟ�'<����A��ʱب��*�m�~���qz�y
��%��Y�R����"�B,Sn�ZՐ�Xҹ�D]aR���͊��:�_cȍ�s��W��5>�G�+b�h�'�Q�gq������v��!� ��?"�LLg�~�C��O�5Hn�F4G�i#A>��X��s�A�f�������H�!���~�9x�[���={6�G��2��r�I,��]�ڡ�J�ȴ�g?�Y\��������fu�J!��ح2<��T;��q8��v� �4;3��
9 �L���©��&�����׆;7��׾r�^0���Ƨ��SM|e��(B��G~����\��wź�UMQ9�,��	��6Ÿ��E%GV��U(	��2ţ(�;wlBk�6��zl��n�� �S�����ᅿv\�(Z�%Gk�`��H��SSSG���V��^A��v�: �D�)=��� ���X6��Wr��䓟���k~w��\Th�E����Ck'�# }'ល��O�9S�����¡��е9NqL��ۉ�:���P9�+2*�+����_w��fkZ���x��Ql��b��9���}Pkl��%ફ�£x>�h�ǜMX~F���dn�U:-��^�?��G�B��)_S�щ��s����6X�B +z���y�,;�e	����O�����Xs�ꈰ4KW��qѹ���������%Í\� 1�Xͭu�.X�W��TN���@�	�C�4��G��hvW.�ԯ'FZET�pi �0v��c�_Lj�ȴ����~R��s�?|�׷	�]Y�����]�� ���I?j�8��5�4�fx!e%:��k�������>|<��'�����Õ�������*w��U����"Sm��Ts"��ߍϊP��L4|	��y0��6$*�&]Y�ǔ��=�d8�,C�h8���0N�/��ึ������K��+~�yY��cbpM�h-���ʮ�m��4���F��6+��:�����E[�k���J����1�!(W}]N�Ĵ�ߗ='r��a��@<��n�y6�]8&te�_�n}�(ߺg��-�5�����(��&�U-VV�z�&F{����J��v0��J�ܠ�*�ipj��q�rj�D�+
l��D����PR�zlGDLۂ~�ų�AO�\���Z���+_�v����U�A�3ϣ�+�׌�`��>�[vs%�!�[u�z��~������7��O�w�d��/���<���1�Q����W��f�b��.yG���u7`���jk���MOa�)Ζ&B�+yI�ڥ��k�7y�H"~O���q�Rڷ>C�B�;f��M����;��ٳA�c�Z�i�8Q��]GW�b���v]s�r�s�N÷��C�lQa�hvO�=i��U����%��佒��~����C�B����u���B"5oU/a�ؤ:@�Gx|�T큲L8X������_�7�.����遟�.�r��VL���V���Gj�uUz�
����V^�q�E[��I��k&�F	enS3�J�=����Z�kaLIf��W�����˗���<�"-qb������i�b260�7��e�T�r������k�ť�x(~'ݭ���G���K� ��?V��e�	Q���G#wK�1M4D��9����'��߷�B��/����ԅ�vaf�z��Ny�6��5�e��� �#rC�;���P�� 8v�C&<6nj^�a����q�RBS�#�P��Ʊv���Yl����/��.��C�-�}��a	rd�� %�*�rKN�
�:T���	��S���uo}����@�ܢF0��T�r��T�
7���Ϗ�j]t�3�D3�L��4�n5,?prV���=�N�3�\�	L��iL�X���`���5�̯}�B���i�a��(߻�?~���_���k��!q��(M��f�{Y>ծ��ط <�g��e1ІU_�k|%�Kp)J`�������4��zJ�{����	���7���"�G̘D5�S���D�&=Z�a�QK�ԕ�e��!��߲��������[���������]�e�Y�%-f��n�[��;$첋��Bޗd�v��T&���/�G�����d�ғN��=뻡l�R�"��|��/�%�_��(ƅ���:��`Y��XV��h���k5,f�i�$.�]q�Ȕ~���.6o9�����َ>�����=��.6������o�lR��_��P��U*H}dB�v��`�ⓞ�Bl}�Oc�3ppd�ܲ�D���(���D�f6nV���?Q�梫��̳X�!3�r<uʌ�
�̕GM,�����S99�yX�s ���.���������蒋A����L �/ڍ��QhB���EW��NV�yB�=�]NF�2�����T��E�lۿ����E����^�
��߾NT�����5厐P�C�^�2�z�"�*����"�k�	��?~����#��Jt��R[�PQU�м���G��J�<�����\��G/:y�*K	�(���,�3�0�w��OL��o�t�����b|�w��=J�F��4����"p@��2� d�l�$V	eg���S�5Е�Ui:ɚX�����¹|&(j��/gI��P� �Bԧ6���,pѣ�����7_������YNR�{hb�c1,k>#��g�Q��[�x՛ޅ���7�G��=�OCM�)�$�C�Pu��G��k�,��KAT-X3�P�@�GvnnN4ƒv���ڼĎi /�]�6
ׂ��\�(C�c��p?���v����+��
�R,�Z-h�hX�j-��<`����$b"PRa� �I�"Z�0S�bkD0Y�^���/�S|�u���7_���b�T!b�E��}>4�j��V�/�O^�B�����|����H��1�V����u�@���ص��%䑙"&W��sG:�l�����w{%��6�T�v�T�5V�?����S���:�#��*�\w��!;���Fy�l�CY�Ly���RO�>1���� �Zؤ���#�Fz4�!Y1��.ϡ�
Nc�1:�Q��Hda�"�ڎ��<�E������az7��m��������z��
�ۋ����%������`�9x�o���v��IQ��E"�X�A�K�lP���!�C8��*��`Q!�蛲��Fg]�����P���nʤ��\��{�Ur������Z��f�20��&� ϱ�aB;첱<)�	�յ�-TV�*'k�7.u�|F�?��~���)=;ϊ)<���ɉ�]��F0�"�T��dd�!�HH΅��`���~?�x�q6�x�ȿ�7�x6�����`�i�7ƕZQ,�o]{>��k�;��
8l��p�C�{S{5Y���w_c8�g%܂�Q�Z���"涊��xdvI���'ی�,q���B&�R�,,P�ƐH�]�j!�Ո(�#��ȵ8�e`l6��']��+��8�.�RXUKк�X�ьR���Ri�j��-�"gdC�}�mŰ����k탇(�G�4S�E�eYZ�f����[ο[K��;o����x�k� 3*������Q��坿o����z��6Av�p㐣�	�F�11���L�3�9��xt�8��!c4g��8A\ Q@Y�fiZ��n���������<��}�{o�UTwu���)�����}��>�������Y�S6�$��'7?�=[�Q��n<��@�V���[�K�#:�����X�.:��U��W��V��Z3]y�����r�)1L�}��F�y�ݻ��k���UW����/)x��d�u%�-�j2�8�/�����m|��FB�C��O���9'r+�Я��gj�;�뱃���	����b�1�������/����1�-��Y��Q���*�l<��߉���S����ִ�҅�ƙo�0���7/�Щf�hh�X�s� �tUL=�#D�n��C�
9@SعR�8eۖ�"�g+�
n����_Q��9����&6]'A�-i`�QIٜ�1�K VYr���L�1m�&Y����O�"�%Gp��,�
���|�T��b�`"<���B1�y��@|!�V��vӱ-����V򒁉 koK�MOs1e2�`GC����K��d�S-R���S�qj����s_KۏW���r��Z��o�a/6�� �<wi~'��71����<�M"��
�JϤ-=�>#�v׫"m�X���|7#Y N���,�(�\-}n���	�DcV�R�`�Lf-�r>5��٘E�O�3SYe�FE[�C~r`���,�?�h�\�˼2�fc��v�1e��z��(J�J�kk�P,Y~�,���
�;��{�4)��/�5��cU�2����b��yM�Z�G�{���C�X�Q7%�.������l��-C�kj�=�^�L-h�-�b�pS��4NҾ5���e^��⏃���1m�8�������tn�
�1�.?,(>�5�S�ȹ_�M`��g;yߴ������b����l
�1Q�߬%cA�e�kMy�Ai�vD&�cx�J��-Y�mtd�X"I�E���x9C���&Β�OC�g��
Lr�q��5�{�հ� bh~	5b�,����H����	Ѧ���b%�ܻm9_O���!d��@��Bƒ�J�f69Y��U�4�
�K$Mc�6-�+��s�֢�U��6���t}�7ѥ�S^�d�X�}�z�6`�َ�	L5yv������\�/;�b����-up��r3������	�Y���B*JS������#!MS?��%�Li:����3iS��&Qm�jV���B�3�vC��3JF�A�p�k�.���h�c�v�L�u��%�,�����T��!&@�31O�l;��a�)�.�>ĝ�:jrjU7��e�l���� 7���+��a���o�
8�*��9G�A�RR�����rt'J{���MN�5��d�#6�ݜ��\a�d�D,�oX��;&I���3g���|>Y ����b�R�W�ТN���|[A�V
d��V�Հ[�+���u�Z2�Cc��:-(�؆�^j�����P3ju7;��6�u��!�ԄWC3a7A���0y�s��	U�0�N2�EExZ�s�����v�VdbҮuqX�{E�|�oh ��CՕp�	&5Q�X��e�f~��U'��z���`
����C�,��g:� �5���{�&��Ս�5��&,bm�h��h%�*)lH߰r��]���\�G��y�ͭ.�\��:�x*�sZO��vsm�@�+j���� �3ϓ�|8�Ψ�E=Nlu��mi��,�ew�|Q����r�)�A�W���%	��+'���k�Y1���]��
=�]�MPP�2�'���H�$���Eiw�Ԃ>hT3	�e7Α]X~f"�f��R
;���H�K^`��.��EK�ƒo��d�99*f��
�Ŭd����&���S-~f��XJ��)�f���Z(����y�٘yNgi��&��{�\ܥ�%	'��_|����ر��^)h;�o�P ITS"�Q��Nd�+MA�X$���b�,xWI��]C&� ����6�����{p��g��֨��/U�5�s���3�����q�a �-v�)}c��5_S;#*�}^4aQi��鉐6Zu�Dk����h���B��<�>��M��T���+rltŪ1����QI@�YO�H�S�/yH�eX�wԖgU$�<��;������d־�\��W�c�J�N�&bKw#���^8�5XV��yY��� �cS��P.�B4B�1d�\�2�RK��I��GP7Mz;�#���G���xg��4���Y*:&�T�B��&})���,'�MY�xj�b����x�ٽ���T��^�Xhf��d磂h���aW��]��y�0��F�#��"�%����a��5Q�IꚲG򋤖��H�%	wD�1������W��b�T[y_"��Si��B���٢���!C��G�g���*ʎ���F�HSi�S���MZ>(����ڬ&_�\6�c֓�4�'GFsF�rX^'�$bW[����N�7�7}�أ�:T.�Y�5	.)��/��7ɸ/bkfy��!,V"ylcnF����kI��`;09n�r�����,(�ʂ��y4��-WV��/��r�䰜"ir`����,�.��9&�����Z_�h2L�6z�&�`��;��P����U1�`��VPk����#aH!''psr�+^ ���9���rbB7gw��U��;6�QW��ب��j��ۗy!CEu�T�33"�r֋�*��k��&����햇ju\ k���1�����/�!y��'�]��T�sZ]y���VQ��\��}�w=fL�[az9Vrh�Mc�%��ИhCu����(:��%���"��u?0AE�x&�M��=���:�
9N�{p��c8�����0|�i���-���<�\l}�)1	c�h�݁sљز�Q�|�|P	�e2j��a��2���� ���5�#��k
�a{W0E�1"��W���k�И�����ĝ�������Gy[f"�ΎB�w�F����ry�蔕(��("X�>���{��`���t��L�,)�;1ʲ�W!��Ƿ�<6!�{��?N<q��.��8�����W����/���-pE �����q�Y���'�C�<���"L�\ds8�2R?Y��XL]����"���)z=�eQ����L�8��g��W����gw��t
.�����(�[������_(��)yE=���k���k��O\��\v��j���D��t��Gb�Ƚ�2��;d�����k�;	����������F���������^�w��7��~��r�;X7���{���{p�+���W��ct����+�a�N��f�&Wk3�~�p��+RS�없Dc4�r���~u�����K��{o�[�r%���3����%B��޻Lͅ��!���YGs��5o&��o
�'��ʳOö;͙��a	#u��h�Q&�TZѶ��M�1ˡkhG�J�d��1���P|����ӂ��������o_{>���?Fm�p�ӣ�n�S!�>4����?˱*��=�c�����m?��-�&&�+�1�u~م�}Er��D[��;�߀��0���"�I�"��B��.������L�;��s��-�:�����!f��{�O�Dy���ˏ�	�굸�~w�8(J�!|����g&����v\��w���l�	ڙ¥g��~�;�\p��w��ߠ��l��s��1��k~�
����}��(.��;V1G���.$QgqGփ`��M�D��y�u�Ȅ5j5��qf�8|j��ȏ��^DZO<��%��wn����>Q��h$f��\��	/74�6[CT}�+���(&6���^3��*:/Ml+q�����σ(����+O��:'���~��9�:���ߎO|�2|��7�L5߸ �07ׄ@̱6u|��:�k�|�F\��Y�M}b�E�g���$��Π$�xσ��o��ٯ�ת�������w���;n=�Qǋ(�R4���U��tF'��\���rΠ�Bn�Q��:/�����]w����β���׏�=덣�W�O㸕�䬔�#��[�S<���8���_�"�H���-y�zm�6[*!����ΐ�jc�R0)�ֵ�v�Gan���D_�,�˱t��S��xIP�`���q�
�:���߉�U���Wn�����������D�4�z�E�4��T�ڢ��N�Pm�ͅI0I�&���#|5<�Z�Q����������.y5zH �h��a`�����ȕjJ�ҳYKIN�Ǟކ�_�U���7q�2fĢ��E^/i8N|�\���,����<�� ���y6�����j;vlǘ�m�=M4��q�ƺNǴ!�ã&�W^7gń��l����<*��J�*�OU�擺Y�p���73!]��O`V���Ę�B�%���7ނ�Gc���R�c����0Z^�����߻_���`ƟϠ]$O$�Q�+�=L�މ�+����4�W�*���FPA^ݖuuOn�!��\��a�9����w��:��ΚXh���v����ג�[y�Xe9L���E`b:��RQcIGb,�%Nn=��X���[(���"�ڻ�ֹ8�k�u�n��|5pꩯŽ��BvbGk'�]�m[6c�3L��p��ER��KLy��Zr���u�8�4tF?���X�UJ����b�ú��bӶ]芠޽���J���VKZ%����v��ǛE��
8&&�"���|^�g�h�����q�[~�ݹ˦��"u�%=6@��v~35������;��4�7=���j5yt��wc�Np�l-��gZTc���o^��7�{����X�Z0�Zq�H�\��xP_�Xr�Ĵ��m�,��a�7%�r<&f�f��L�?�p���l3�Yg�ؽ��!^�oz��}'`�ګ�G,�+.��>�"�>|9N���e�0GrX�k�i����Z�ZH��t�n	���؃�}�
��0�v�Jƕ>�NΥ�	f�9Y����u_��?��I&�g9�¹��A]>�����o�����;Q�2b�#u�G�֘�1+G�H\�T��b~7�|>��_·nK46N
��]�㲋�����n��j/��W��y�w��O\���x+yR4�tξw��\���%\�\�Șah
�֓��6BKH�J�,z�����|6?��y��V��A�����<��^��?݅��;kN�㺯��]�?
�z�L�|� �;�߅�b�TG&ЊM!�U��N
�ɍd�c|r~p�#��&�]y�&��]�ɗ��^�-�o����L 	J(M��O}�Q�Ys<vEں{�z�$������	<��^�i��V�1���em��h��h����Mw��-<���P[G�-�?���pʩ'�7 ��~��=�1���?�c�uڙ8���`/1oxRۓ�z~+J�1,�^X�8�Y)_�c�0�����J�7[������U�}���Ҡ
�6nA�H�}�I��ûerD]�{<Y�T&��z�V�{�"Z"��<}�����N�yL2-�X�t#Gf����t�FmǊC��ZA��06=�F�m���y��&�{�!�6b�����>�r�iN4LՕ'
0���P��N/��61���c��0��Ąn������ڔ7j��ʽtEM<�m/���S�L!V�	�� (O`J��]?} w���L;�ȊI89G�[���s�a�B�n��b���J=�.*�5��07�f�&�Lݣ�95I������SutR��YdS��Y���4�b�QlZy���8x�X]�ZH�E����f�V��� M�_!3�=�Ֆ�ntM9�b`�R����{O���k�e�6�aƕ��[BI*5yF�¸��W�8��mkg$Zn�$���wCK��_�Gb�n�BQ*�I6�6�r~(����n�����8>����2Bȸ���TC�j�m���fՙ,�/�P�%��[��$Yu_A$���j��9e5z��:���lƒ��<p0�O�g���fFj}v�����hn�>r�os:L�j ,�,#�VEw~���S7�8��s1XRijK�L��.��[(��+�6���8�9I��+Ô�P����@��*�дgBNfڇ�R*[�]	�ѫ+IM	�YN��k�H̸dȘD��A�f�w`��v;�?D&}/���6|�,1]1m+%��wuA�W��>��,:� �.�9r%���P��"*xn�/0ĲH�%�i����3YעB���1�"_Y/X�i-ñ���Nb�gW+�px4:ME:i��r�C�%�]�ˑR�g����4-k�|6���AH�� MFnv����L'1�_o5ܒ�0^��q�E�1̙��>����%�D X�����m,??���n�G1/��4�5��}�}���[��(�=���0��~ـ����I�Ք:h�<jXGܙ��_�N��=�S=6`cv�y>���{�s�[�����g�M���Y�L�C���Z�GuxT3��-:bAl�n4�I�T��w�ƈzi�� 2ZG�3FA�^]�����_Y#k_���Y��K��Bh�E%�d�%˲���~��k����U�@�ڲh�bT��G2�)CLb;�?��ɩŶ�,�~i<3V���|��	5�[�N��~��:�X <2��,\ʉ�x2��vD>�P�F<��M��^̳F��l�'X�7�XԀ�G��K��YMg��؆S3�dwT�t���|�������}��2{� ��^��J�wy�PALu&�v�Y��ǒ��,�a�t��J�����f�h��ҋ�9�\D3��i󖬒l@�M�`
۪UK����/�ݬ�Yi��l�T�~��lz��m:T�k5�,�\�[�[�i�X�	��y�ġD��L_��L&��TL��M��fǓ&A��ep=��\7�f��$j7�a�Sd�Q�PP�D$$E�m���C����󥏃���1�ť���c֏r"S�?���5�f[i�>;0˫c��E���O��n�8����3� K��h�2��Dq����[�J3h��.8Øb߮:�l����P��hE[�0Ɏ��T���5�A0�\�J~_Mc3����J*3�=����Ũ�v���Psj�\�T�Y'jj��tvvZ��e�Y�+�0$p��.c,�����݁ߘ���R�BFJ�M�S��I-m�vc��u��j�|l�8��i�]*U�7baP�n�,VÑ]W�(��:äh�h'�����I\[39�HLN��&GՋ\<ϵ)�L��h���	]�^�B�ߑ���g����#U$Z����=�1C��Sj�����g�7�I=F/����� s5us�����"�֎��쎒PkRY�C"�?��ۊ�]m�j&��x��<�Y�K�+:U���k�t��f�f��,C��5���c�%L�%���Tr�^ʤ�G'He����v��R{�� c#Qqj��z��w��ۨ�b�G�I7����`�E��8�'aI(�t�~�i����1��uy�jf�.���jO[f�����D�܍Z�wш�9����~Cch�]��fn�5�Pt�&�DU{����/�FzS�jo_�s�xz��tP��Ư�g�!���j��p��?�-O>e�J���e�%�ݘ�1��4�3�d���Z��\DzL2�~���$��a�Y\��s�n|�~�j�l��Ŗ���0��B�%�ϬtP�{te�eT^�bM(ܱS�����SN�\'���$J�1l+δۄ��4=]t���B��	�X�UC,&��f{�+VL`�ʕ(TC%Jcy`�e"������ڂ9���V�1��;�Be���W��>
f���n��L�g�Zt�E�C�d��I�Z�Ƥ��zH��q��VKwp�
�U{f"�l�TK��0u{�ڤ�1j��hʢT��-|25nd-�)��U��wH��1?0�5��G�O�n��<׀�N�!ɉ��P��R!w�[�$�J���!��APNv����Z�S��	v*��FC�ZM�����[��<l�!A�K#�9,<��A�M�7Z���o��p�f�W�>��
Z�϶��rrg ��)=�CH��}�J�{B��s��'iڗM�jm>�(�M��e掺I���	��YE���ؚ٬՞�<K|;}W׿�wA�"��Ts�m�=ǦO:�ݲ���B�S��jwǦ⩊�S� �-��p,ڎ`�PS���L*;�\Em}v,�r����N��_�l�Z� �g������ɤ�ϜI�`�g�zb,&�Ȗ���v���G2�ˬ�h@S��3<���1�*Y2S�Q�iE΀X��Ƭ�����hu{~�Á2<o!�J�@��]���=�6�<ƞɈlNbx*L�(GU)���Sx�hV��v_���a�}��n���ps�0K%����K�kL>�)2��*�%bIP�źP>V���׷�%��d�Y}��\���U.>���YI���j5EӸ�T�U�`9fU~��'8i��4ѡ5e��quc��D���$Y�Q��f����4�~^F=f�˘m� ��1�	���`Ǟ��9L�U�]M��,SW�)m`�bH�*�}z��2�s�d8����KQ|��U��٨��R�\*��@�VIg�"���)���xP&Z�`�I�Q�X޳���S�@��ݘ�������A��C�=�m:��i�����g]�f$ڔt�8gI�.�(a�gԣht���he(��j
z��,S����������ʨ'��MicS�d"Q���A1fيI�P��pkʱY��H�-dHk"�Qά���f�i�bF{e�:�b�ٽ����1��Z���O~.��mHfg�b��"[7c�.R4t�PvB�S���gFN,���4��FMP&�K
��{��4r�u��{�9�t�qfy}qT�gO�56|����~g>�g�����=���
��bQn�>�@�'�t�5�fo6��o�Y�)�\s�k�m�d ��G��f )`B���S���ȏ
���=�B��i��a"�@�0--w)IV�jg��0��3-4Km�je=B���d^[	Oש�B�u�NS�V��
Y]�$0�����ޖ����2�$0:r#�Ly��b�fy���p�H�e=�M��3t�Y� �D6Dq��
�m�HyRR�Fj�����ܘV�i�΁����P�ˏ��t�m	�����)���!i�l9H��OTS�-�Z����I���+5�:cΣ�.Q�����NK&�.�2��_��+�{�pjd��[��\�<fe#EE>��06���רFI��@vl��x~>�D }8�y>'���b�_������J_�fTE ���$,������Q]�mnik�x5�g�@ǩjL�����S�F�l�+j�԰�e~�����*�[Q���\D�*������{�pN�4�:ن<��X��.�U��@,'1��b�9%�˫А��jH�|�Y�c���g��� G��`��t3�4_�$�4�i�D3M�}%�=��E�@D�1fs�����	ztݢ��rSC���RfB�D d��_�
x�����j�tt�o��;��m,]o>6�GY����x,�NytT�挋5|m���pJU�Ϻ�cȻ��E�p�Eb%lD�Qv�f;%��2�8�o)��9���N�xEF6Mb:�XFY�܀����9;���Q��M8$J���&|��;�"��l�*�\���Z~�d��d�A���1�;����_�����j]�p.��e,'����Q��I�I���D)[)�4/�-:2�,��r�Y"V���7,s"�*�zu���� 8���u%{N�k�
�d��'M�O��f&����۠)Hb�VB�9�T�ihW�*h�A�(���ޥ֘�?���$�+0�6!/!���`w欦�65�ɓ�yyͼɵ�^(�/C*|Ij2�� d���u���NL��TK�r��Ӂl$�.�3���0f�%�R�JD�%���s0&���G`�,��؀%�z&3o#G�5�-�:(��+g��/+/k/�'�0ǡ(�f^�C����k�(w=8��7�'��Kר��-��p�Zu+k��t"s�U��O�AG@n>ߑ�5���"��vC��	��0A&(1�SqR�������f��O6�Y�T�+�u���ԛ@�SG�K����䞺ih�H�^W⩮�0W혓�(X�A���`�.8�RDCE6M�`�]�-^�G�rd:6�L�w�ɵ檓�I2_ej�2�s�r�5��h�S+�y*0C��ɤ���b��b��Uu�%a����[�=E�u�[�9����u c8j���cCs4���|�/��#�8$d�]4SB����=�;m�}B�{�N�i�`�+���Hh8��	4��8�<�иè�e�ш-���X7��	-'�̙�Yģ�ڋͳK��Ԉ�蘒��`Q�}���ibx�X	mG1	���E^o���3�Q�T:�}��"['��,�����Q�nhh��:�M�I@�fV�(��\��ȘoZ��(�{��q]ߓ#�����6�v����5�FNO(H����b���z"���Wa$ECО��B�]��X)��2�<�ג�9����O3�f7҉ɸS=]k"g�+M���?��S��(3a$Z����d�b����	f{�q'	�'uc�IO��H9@�U���J��.`d	�����O�V&b1@�s�`tc�\7�ϹCb�9i�T�Փ�CS�x�ߡh��Wn^�"Q��y?�Ė/jy�Q��p�-TGdG5v��D���f�i�b�;���9Vx�DF!���5NJDǸߍ��|�:��sI.g�.�0B��F��]Y�Ey�1�gŁ��j<�q��0����h��>�h̲mu�K�����{�%��A�a��e��1���T�݊�ĵj��YBN{'	،v� 	��ߗ�):�޿c��C���׼t^��r<G= ����~�|�=��m�[��"�yG�۠�.�Fԏga �!���W=��:k��� ��Ҵi�E�p.�̟x�BŐ��ۋ�ʊ������H� I㚝h�b#�^'�B��=O��@OuQҸ�=H��5�����������S�v����Ǣt
�>Wұ�fKE��g�G=���C��Tk0�<���v|�ǳ�Ug|��z�0�[q���\vT>�|Of�4~��|+V3��h1�Ӗ�Ԛ����
�o�ƻ7�MC�9\ks3N�&?��������a�El�LD����az�?�隴��/��;�FF�l6���O����?�p]o�k;w<�X�Vav��7O�����-��M���շ�cc��x�ٍ#pm���6�s�|�������_L��%�\	�\��_�η�������������߽`>Ƶ���^��7,w�,������۱�T������9�\p�,�а��r���߿�'����ј]h+���^�����6��f�v}����N��/�(�l�Y�c9��P�0�(��8��_��:Ђ�a�S]�k�A9�ꄫ
��rX��2/?����A��D�B�GqS����Ǳ��)�1Q��e�x��I	,B�l�Q����c�ޘ(V�rf7��/F6��wʬ���֬Amz�����n{E��n�y��W�57s<�q�K�D�^�Hշ��q�qL	F�T^YL;�3�U2����ɏ_��|w(_*�_��bg�b�8�4ʗ
y��d�/�(�cJ0:����8��b���0q\vC�>�sD�'�v$ʣ�>����e{�cJ0d��O��xK'�\�p�z��ue�JQ��'ը��7��q�	�<��4M�M0r�eJ���/����a��A��˭��֣z�k�����Gl$��KO�^�؟�`���8�#]47�aG{.�0KGq�ɘ7D�� ?�C�����R1����O?�`��w�r.�����V����hjO�G���ڗ��Xf�8��_�c �l� ;vY����L	�Qǔ`�_i����r^�c�1��U20����5�����܂1o-^��c�s}�Dq/}$Ird,|��_��1O0�Y��s]�h/����e�d`̋O,��V�����Q�,�bj�Ʋ�ǔ`d~Vl��5�?D�Aļ&��I��|�M������Q���.'���(��m3�	�V����jy�Ϝ#��.�qL	F�[fa��o��,H��lCCCڈ��l.[ȟ�����5���pS�Q(��Z�P4E�NҞ庶��z��Uv�zY��-��2��cC�,��]�V��Qǔ`\|�ş���V��eq��1{�r]���/���۷�#BY��7��n,���K�X���T�3r�8���6�o����q�eU���8Jc�ڵO�ǔ`d�h��c��W���3j�    IEND�B`�PK   7��X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   7��X`$} [ /   images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.png켉;��?\_ϣzR�'B�OE"b,-�����f�v��Rc�Z�P#$��R�l��3�c�Ⱦ������{����}_׹|���9���������u��;v�Ӿ
7ܱco	�{77��'���������O��X�y���[�;D>��wV;�0�Bk�D�ۡ1V^�;0�YG7g�����Yw/�D���;��І_�����D����,.����? ��?v�@ў=r���>?Ot�8���g�8�Ko��ve{��;��M��g�d��&kܖD<Йpo����k,ѧގH����@5F�G|�X��9�@�j`S.�'��[��ؿ���\�m�݇m�h��Jx۵9w���{�D�c���W��%\[����vn}����ma��������Ƿ}>�cN{��!������	�#�{��.��26��������.��qDSx�v���61H�~���/ڈ���V��|~
t�Kk���!Q츨(��?q6��k>�4�r�K)�TnG� ���*�E�Op�@�]��\�;/˘a�y3D}?��J�������%�����ٌ�<�U�Rb�pT��f�%�\��$S��J�d<�T%6��#AZ���ǻC�zs��0���?Y����z����c�*�9���ޟ(8B}�Uv��K�!���W�DzS�ڿ�¹QFn���\-�-|�&L���X^�M֫�-�d=꼒��t�?�>,�����3�ah�1 Qf��qːY�����)J�	B|U��"����;h�5횇�p���7x��-���"ǵ0�Mø��3j�3��$���6RɟVS ���Y�|䟇e��&m���>.�E�{�.�Hd�Z`����)�E��w��4	����ۦ	h��;���b(��?���3�nԛijiY�7���[�f���ʢ[�M��-o`+��]�S���ḇ)�˨4�`s��ϐ�5��i=ΩX��\��0�żӸ����Kpx��J�e�ztW�J��erC})�� ��s�>��+Ȭ�?'�a_wu޿fg��0�*�{2�as����@ۈ̥/���pK��~p-j��uۖYo*�%H�Ab$rp|�,���6�FX�0��y=�M4n�G�'�s�_�e����>���x�d�k�������f��$�D�����=��_;#�z���c��$w�����O[�&�V�
��?�ݾ��|t���A��U���à�Ϫ^&��A��uص���qX"����
+u&��SJ�V4S8(�}�")�+��i���k�<j�~-�=w����1#��5�E[�ws<7:)e�wmt�U�#g��r�1�jB�{	*C��/Z�X�����V���E�i��Z.���E�pa�L�PS��<���w��C�Q�S޹��G���)!�*u�nˁ7,�o�n���b�:u�J�����f��A��J��'.f����O�-�g��8B��$�PI�7u���;����z�>{V����K|��Zy>A5c�
/g����1�Z)6T��|�/*��,����MD�8֒��9��++�����4�`z�Mک��e}����ќ��CYI���
�Z���ŤTe0-�FY�=8����E�A�]c�uc��^�/#��F�R��kqbi7�jԯW��U1m�/̏��bh�u-m��y���W>-�2�߇	M�H7ڈ�2{N����b%�뜈�M<�S$��r�Ot��e���K2ǯ*�|�í��������'��k�������:��a1�����J�����������&�#�&W�J�(�bUOx�J<v����.��rcqC#ĉ_�E��f|��%�h0L뻸�3a}��a�k��M���<^���~(���`'���"k�	=`��5�����^�o�EjB m��h*��ɡ�{_��'x������R���f�����Zm��f�4i�U^��AT]��!���Q�UZ/E����ÁD�J+��նܰʶL�%H~�;�g��ƢGF�L?�����ť}����ōϦ��?ʱ�c�����d���^������k�i���IL��@�dh27N(��ԿaUJcmm�O��y�w=,0OL�G
��;~|�*��Kc4��M�7n��`�c\�����g���Q���I��Jg|f���v��h���)�՚���mr�)N5ڤ0�e�X}���{Xm��_�ƺ�"��%�#ǚ�a:��$m��ŗa8�$����N�B�z`���|
��q�~���A����ӻ=jić�Q}{s��6[�
o�J�$���j}�~��P�p54�!�3���A���F}�©��S��C���q��9]�OPY�v��r�Y�0�gD�0��gLm*+�`����pS�lp�����I�2�rP	~!�̕ߔE�<F	n�g��a
L�)ݽn��}����B+	e�h�s �u�L�j���n�t<,�M6S������-�2_��+@�p4�Lʾx��^����p�U���q��ҁ�}!��Ya�� �Q� ��ʪ�S�oC������������l��Okx����m����V��S}<A�mH�\���E�ֿ-j0D�:�̼Lڸxh������e�T����Zl�\7�I��n~�b77�N5i?[�SlD���6��$�pJ)�>x�ܰ6�:�v��!�	��J�"fz)QÿbJ��@��N[��niI�jZ�N`!=>��#o-(�W��\�:Β���	�9�qyӒ-t��4��v4p+��a�7/yF�0�#�j�;#�@�_2���q�B�J�Be�p��?4��j��n*�����3_����j���*�~��v���7���m5�i�!�P�V������P7����;~�M~�2=W�q6RkP��*��Z�>r�&Xryk5,�6�qJ�ϖuԎD�z�K��򥹇�+|�XP������HY_�(�X�ԭC�Λ���B0�������c��f�M,;RP����vQ儅�&Z aa���7��F�r�=�Qu;�HN����a���6��2�\��,Iq�5ăj\���n�OPa��)_Ɏ^P?���Iл�CS�� ��n��M��f�F�AJ�Q�jhȢ���1?P(i!2��"Цx
�?��iAH���I�8���5�Y ��a�|�ƽ�O�:�5@;`2,�1.&�M�hh�_��ӿ>� ="	�I�#s��ʝ����������k[���ͮ����ɗ��Y��6(�_+Ps�zuW���k�y���H�'�v�����wN�z�7���5�5����ˬ˰I@�X��&˿G�(�4�0f%��O�#�e1���
G�3�w�8fU�Y�k�g�6��M��m4��'��L����*�G�F��|]��ߘ./�t8�:oYԾ_�`uRRleŋQec|2�=��W0����<&��"��t��I�؍�6>tk�����R�|�U���񧒣a֝�,�^���>_jo�͒��7�� ` :OiI����X�C��|�_>�$��$Ptl R/��л?=�;��g��*��5�
�UN�s(��w�*Ս��ΟU@����+��*G��)���Y�x��%vUލ�X�uS�"X�#'P�O��y�_�r6JB��7x�~b+�)⑰��&�G��[K���ק
f�<�'��N��y.R,�$bΧ��ʬ�o|�:�g`�v�
s�	 �wp��e���r6�Z<�	��34U�_/��2z:rl҉�F�ޗ0IAkv�̯a?�r�b�g@����i�	�j�N�N�?M���_��I�I�KD`Re����3�z���T�����H�@���
���i��G���������z"q���Hni��}�Z�G
�,��)[�=Vi*�W�Oc�*�j.����t.�V���,�t�a��
!7S������䕘�ƨ�5d��uX���y�]Tpd��LgA���`�:xgh Wm��n���g��kȹh������QX��+�I���a�kډg�z0���n-�Xډ��xOh���b��Sa�iz���s}�������l���8X�ZX�}u�<�mpT��监�w\p�Mi>��=R��I�R0��J"U�0,+ng��IT�FG���C��ɭi�i��%���r�9��\���
Ǧ�-<Ş���C}�~����f��|#@v%cBLS�� ��[P�����;� c��=���QS��_|ɓ"��A8��6H��X�^QH��t2�nn��װ��gp�V��Ν�<qh�J� O��FIH�T�<	6�`^-(X����v��V��>�����%�;K��Ò��t7w�DPn��[��ZF�[_�8�������H�\���ݘ��0�`ב x>�[�\�⸓�i���Q@#�C4���7Pk#x����F(	�/r��X�����ɽ���D�j�| ��k �z���c�$������yiܸzE",����h�C�����b�b���D*��.�������[]��\��]ӆӊ�{V�VN��0���5k�$��Ha~��s�ﬗ�ޘϐeW���r� 9}����f��i�vn�:T��in�R[kq��	�1i�|����ˤTN�O��U{u�!{A����w:���l�դ~LҒ��\�� }�!��|\�I��Y���$/�v���ԓ'O�񰱼��kK�Z7�H�W��$���G"�0B���]"Gg�ċ]�.X�;n��6R�{��Q�۬p����G�'��f��6�:�w-��@��>�)iii`m%�^$�\��Bx���I�ŉ�xE�������N����œ�h	�+�>�uJ��D�0�@�}�����]��}ݣ�k����%�A�5j�nq�oY�\��a��Z�8EE�q��u��E͚ C�TV���Y�S�҇'�I�,V$�2[�E:M�my�D&?7T�A#���;�� ����5E&���4����,�;�4�e��̦��
0��,2�v�|���ŕ(6,
��s0�E.�Ҡ�IX_'����9:1U1"[�ն5�;���_��R���u	�F;��uQA��������b��L�'�u�'^�����J�ƀ	se��?E럼!�>���r-�5E�]��h*���!��i�#4�ҟ%������YS����J$�=���'�L�Ȯ���SƏ�
��/.M>}��\��+nll��3�,�=<~�b}u�G�Z.}��0�}" �ɹU]vʹ&�����S�FK�<4���'�]�xXZ`�T��_4��sW�b�VE�2`�b�88{	�T�AS ��Q�����,�g�䔟ck�m��e���P�
m�.��|Gn�Cٰ���TTֈX_��"��'��"JӼ0�a�{25���6�Ȩ�_�2S�k�m4V�[[$c�� �[j�)�m��q���R�,�R��D.�.%{��b"��ݵc�M��_GiJv�j3`}Ȭ�s�T���ӮMz�wԏH�O���7�R�Jt���F"M4k^���b-��5�y�fk)?��Ł
y	��x�{:��V<�r��	�5�>�o�fH�T�H��^6i|{3�,�ɞ�CV����c�T�e�8a�c��d�>��Oi�.�9��=��d�Xt8ȫ	@��a����j��H����z�.`������!�Ҙ}��U�E�1�zfY$3��Ėё�Ƀq���#�'��@��I$��d�Lk�����`R<M	6�<R*�z�7��x���jM�iv�my�?���,�nJ{��Mk��|��0{�����4@�@M�8�������[/��Q_�~-�c�ӄ���OeB<�Y)�O��ǉ%��q�L$�)7�)�hm`��Hz�
�Z��#�/�g�zc�{=�B5k`Pky�ѡ i\߉8�t<��0 6|�G����s�X���E:�$8n//��Z�A��;�� $��Q�؊t�� �Y.�bk71��K��s$��#�s�A������W0����by���vS���.P�ό��~ rK�$RJ����C��e��\:�d��W-�r� $7��R��,��(.���re4�:.N�g��g� ΍��{����!޾�99��($f�Xl?j�Z�LR�t�m5�2��gk�ɗ?g��DJ�1 �Km�ȅ��j=.
�C�$�Q���z��m�C��b�a���D���T��)9�ڇ���Aޢȩ���� �b��B�s�髬G#>��ֽb-��1_�)fw��"�G���K7�< 5݊�-��6K/A���.�*�kTK2t�������K��W��Q^�@D;�L744d�dך���� {�B�$RH]�5���Q�cw�k1wP/��}̦l��Y7��� �!���.wAaasd��~�܉���5���Z�p19܄�������ȟ���Q�xc�����Ea�A!����-��3��r:2�}:B�O�p�qz� `\�Gр���TTk�Q|�N���E�e��j��}�#x���� =s�q�R2���	��!��w�:����#�y���Km��	;�/�a e�l��J�-�6[w̖�#�.�H�Bb̫^��gO��Y�PX�o����<�dl�������igC��` ���6�Y���"��{�7dz�K�GtN�ⰦR �w�R.�-<68s+fC��Bv����Q(@��_�re����}�kG{-^#μ�����9�Ug��y��I����B�����6���.@}��R�J����&��L��T�$�Te3o?����H�c�7�ˎ�v��թ���ї��кHd�FM(�� N:���_T΁���l_~�(�8�\KW"��H���D����l{:&S��pǾY�8���xq�}�P ��i�E1Щw���,��
��O�H�D��k1��V�`JN[�ً?�t�9T B�.�4=̃u�e~�G��u��	��'�Q�F�4�h�$�5��H�q���	��%�Z��g���u	V$�o�i�ȶ������ɔm`�D�����)��Пѕm���H���t2 �q����r�N��K�������=�BI�E�"�Ͳ�ȨPU�yՠ�i$RN��	@���j��h�yS9��~�b-�x��}���Z�J�ċ�ۦ��K��/N�3M/_��,�,X��',�dh�͏�}���[�@m���\�a�Sah�����{q���ĜQ���]��+�	 ��H��E����H+P��L|d$`��keJ��P�F�s�`ˇ�-��gP��t����\���R�>d:�9U ���Y����ר�N*�������A3���� _Aw+��0�FE�Ww1�r-���)է��2�E�M�/Lrn/�I� D�~���d�"+�ާ_���Қ�w��
A+��i�wI4Bd*��e�?^01���!�B?���P���X�B�� \����#�&��4qh�������,Yy��/qQ����k#o���[l��=�c������zY@��W��=b��~��b�`�L���'���v*\��C,X��-$�!!�/����?��K�wp� �R�kj"l����-ҹ7�f�A�(�%�#���6	_^��5��f�k��ɴ��s]�	�%�_�;��Ҍ�� �1��:s!�Ν;άe&Y�e��L����$����������9'b|���+�}�)	��ሺ8T��rnn��d�
<��)�e�h��|�	��G�}c?����]���Z�<��ZZ����\)5;��\��K�%$�4�����\���i�(`� �ce���0\)�I� ����?�gs�Y/��T?��j�F+EQn�۵�Ҏ�E��ac�g�Y#��b���Zkw�_/]��*
h���S� l�Dأ�<v��Nv`Kd�_W%��y���f�d?c�\]YI� #�^	����-K�av��K�B��p��-�_������-X�/Tm	� �)`�|66�&^@�����,T����G��2/���{�����ۥ3��W������Ȋ��[$�w�#s:���Z٨(�7�P"��w�~�n���A]�BY��sB��F��럺%{�h�P���p!��!��v�����8EY��nd[�.�
�z�4`���HDa���fw��e�L�* :�L5�f/���"2�� M��H�o@��D�,=�Ӫ���\���*y+u�p�v�N���CM�q%*���v�E~��M:�"A�b�����@� Ѹ����N�� Ye���"���^
������VL��� ��`K؎�a�K%kNo-���/�����Rs�~�o�v�����3-R�}����0��#��r�i���e�i$��k8����=;<����خ��W+V��>Cd�O�>���\i%ӵ��h��Adk�b>zע���"(��5��T�u��d�f�)~}F4C�#��)"���FsY+$Ҽ˩Э����Ъ�����e5��A�U��'�u�VCj�8��$���[99h U�J�A�,3��0���Z�M��m9�\K�L�]e ��]M7a�?��(J�c<`w�s��T+O�s�^XMi��g��?�S���-��~du��V�$�@�[�9 B�������^��%���H΄���<o��֒,+���~���J�L�U�ݻT,��+���؞��G*����Yv�]ߡ��ɲ�~�tځ���[s��5�j�	73�{�-i�(���P>�[�KMS_K?ӴWѥ�k��矠!��I�Ǳ�7J��8me:���pv
A!��]��2�	M--��C�nB�3K�>/Sai@��=מB��J��I$I�]����9�I�6qi�a��m\�_y]X*yrxC�?�T�$0ӄ��O%m���fAC����G�@Vo�a��gO6�e�Т7�8S)j�|��0��,>�~ z�c��r��k���ɰG�@UHA�b�=���OF�2��=��H7&�Z�"2�$�q�]� �G@0MJ7���]<~�7�teF��P��d.C�Lߘd������+��L����w%X��`�tg���}����L� �n��y��
�
�5���WVn�/����tӗ0O6S�O��9r���w�O���u����A~�2X�j�Gi��Z�(o��7_���D�����w��H��(�$���`��	�6U%�lR��[��T�;�k��-P盇!S��Hm��Y�W�1k�?�M��n�
ǁ}9�6�q)���+MM��2�;õ�y:
v��7� _q�k�'}V�c��,�kV:���]�]�P�_ld��ڽ�5�*6\�d�A�ö�(�"LL��9�F���-�Λ�(�f4�F`�e��^�Q:v/��trm�Y��`�	ɓ���d?���x��S���ט874	�5�]Q�i	��N�A-�R��*����t1a�7]Ry���yo��b�V����Q�1m���i��"B��A��ݾg�u�Ud��	�����pDc���!@�Hn^��_$��<��&��p"��)��(�����5VGZ�I�����A
}gT'����F��11��ͧk�m�N�׫F��4��I`
(&�0?X�Y��`-F�7���?3��n��(���< %�X�Qp�6���mM
܎�D�c�(lCo�}&���9c�ȍĆ�0�Ȩ�='%�eO�{����wf�z��y���î�j�F��&o��x�Z�zMP�6��'��[�w�t�(�BB@2��:�A0�v>;4)�8�H�I�8K�Ȉ�Ol�Ě���:��P�+��Z;$r�K�y��{����8l�6z���cn�~�{5+��`��'`���yo�	\��;\ó�"|��M���sd\�%d�;��~=�L{6eᰋ�x�4��,�����k�DH"�<iR�!�7Nb��;�x�5�s����a��Du��Y�Y&�1d���v����1ZE^��6�;���*��7�}�)v� �?�K1�yw��8gr������n��b_�֠���V��!�{1�ʊ��X��M~0�&˞� �S�;^��t
:O�{	�c�nƍå�y��/qLm< �� D��ôgh;m���V�����g����Z�"���v�ç�eN��D�n�8/�T�/��]K�/���x*� q�C��&:")����!�M�@y}?������G�ث{]�c���H�l�����ɵ������ɈL�)�t�C�+c���.5j��|z\)`���OC������c���+��C��?J�)ʌ�@���]�3�UΓ���o/�O���%���l�E�Ѷp)�,�ɜ��|�_W���'cX�YD�;eG~��Ću�0����0YѺK�s����Ǖ��MesU�QzD\�B��o����	}��1`�;���ՀCBҬw�����U(�ΐڣ�����?��Wǩ�Wkf�[<���C""��@���VN���h�����= ID`x��W�6�8c��{��Բ�;�7�=����LV��&y9��҉
D��YUl�����h~f�jg���~�sU�n�5� "{�a$67Ț�����uU ���7�E��;o'�̹����_}x������e�D�_2G��S���y�÷�[��>����`��n����rN��
w9C�}��9(vH�t�,��V�>NPX*Y� 	��W����XZ=t8�*\=���y�4�G�fu���e� ���5*�Z�Y�tl#\��5d�+Q��/����V��l�`ĸ�{�7lt]I��RU�f~�nտ<��0!Q��<��x�NF��� �ͱW����]�=��k5-������;����'��|L�(�m��p��j�^'������/���Z5Q Y�����=��1�/ꞃ�����{/���s�Ĭ���VDs-������{OZ� �T �vV���2��o�C���6.jj����%�t������XJ)�	�q����?�4����2�$iv�x���X�FxxlN|;M����������F2f�� \E�A���j�-�DI-�^�B��A�����	h*�Y�lx��A��	]�d7����g|�8Ju��rƩ{K"f[���TF���'	�HƓ Ti"�D �,�##���,|���ԛoO����و7-D��&�U���l`�'tt�y��\��A�*�$��]{5�� ���5h��	�"u����"?[��: !D���3�����@�Y)JhU2Su��� J"YHH�g�뷙^��Ei�U\u�F��B�>��ް��F��������j�1P�ғ�ّ�@/ʾ�g�b��>���bN<-
�����e;���S��Mi�,P��8�ͧ��n��ڮ��"Z�IxC�2.;���F��s�Sp�ǹ�i�k��'���y	�3��X�C���W�
���h��3��g��B���s��'슨Eٝ��g�W�T��ˉ"��~���L�,l		���#Z��uIS�Ep�O�������WeP��֤�����F�C�ܬՙ�]*�����e;�껡|G��w�%�S�w�Ş��pǏ��*�1�S�U;���(�����*HT�W5��+h��:�/u��D �M�[���T.A������pϭ�/n��{0(i+zx�>�[�������$��u3�}�q�XT�k4��M}�(�������4{GJ�X���a~o�n�ĎE�3�-�8Ne�j�*�_mg����>p���>(��L3|x-��f`����p!p��+'���N��x�{�M�$�=�~JC��^��4x�l'�/Ϧ^�eԎ���+(1��YQsγ�9�d 9v�*Ψ�A�n�P���8!�1���H����o�P{"�3����<э����޹�7-
a�^����\�;��DJ����E�B�G����;O
��w��FJ,,�~pdR�x�=O�����[� A�T�M�NlB�4e<�S���k�y0�#��+=3F ��)}���Ϛ�a)sNm_�lڑ`�Z�x�-`�/9� �[��l"׫���d��L�Լ��L�U�#�^��5��L��J9��
h'�iij�Ĺݣ$���q��tT���hJ�͡�n�.��ەq�5�Du���Qʭ����ak)�b�
5�y������*�5ۿ�����$Q�c0�P�M���^��.9�r^�����h7DLL,�����=�U�
E)?�i(!g�+p�UF:�oZ���Zp	����7�JˍRhk,T2��D	�mkk� ��oy���������E�c}���aC�d�&���aZ�q1%Эzgؗ���.+�ܩޙ2�{|�����}+Ľ�� Ǯz��q�;`��������zRB%���R�ͯ�r�=���9R�- �^a�o~�j��)͠E&F�/�f>�%�> N܅�_c4��B�"�cajg����-��ph�FʜR�_8�֋��+�:���ޝ�+��FY���qnY|�����=�V�)���;ĳ��+�����_�H/;�,	�￧4����ؿ���D�T�+n�=�W+���F
����=?�d�S<ـ�Fuv�"������Hq@�>g&��^o�Z&�/?���f�%'�Uٱ�e7TԚx?Kb;�+,�j'
����p=��eN�d<�w �S�E���$�Tn��6���J� {R.��Cvˢ�T��=��JXJ�J)u�u*����؛7@ϔ���LKB�J4�Ji?�.'���<`��-�S:j�Q��;NL�ƹ	W��s��WM)eyEC���3��W#y�t�cz�*x��6߃=��Cc�MD���5W�?���8[J�*�@K�˾���0C��Vh�x^��[�s�����p�	"��D�I���K�Q!�s��P6o�w[����3��)./�ͩI�~��cH[ʕ+V	R�>�xjݩ͊��
���dq������;����3t����d���v���8U�ک>�/���`����,�~�?�}������P�	 e$6lo�o	��io��K��H* e&d8R��f#�l�׺d5yn֙�߿��j����U'
���DW6,����SKU�m�'�4��U�`jF{�٬�#ǮJŶZ2KT�(A���r_��KB������o<������V�y$�-�FE@�.<�-��撐���r�Ox��aWZ��&��Gt��L���!U{��t�h����P p��ȡp���_S���#�<��X��e�ƩC�Cf���N8���ܕ3�y����o����a(<<�`5�1������j��>�A��j.�[U?�Ҫ���	��[�[���
��`4
���$�Vl�[4��j�v�ߊ����7m	�D�v�(K	�̻��l�-m��y��R��4)��)�Ӫ4��]�~FW��[7�1��N�8V/�=���Fr���EwP0L�R��R���t?����?�9�Հ��xR�D9�;6"��d̼Z�O�F�&t��q�|�ʵ����Q����`�y�d�ܨ<�+�=�պ����f����.��~ԭ�(4�������z0^�>C�Y�pB��� �����!έ�H�1�{/��h�2+�WX��*
'߃��P���_��}C�Ȉe	�爝 K�ɕ��j�H��!�����/w��l=�˸��&	X��
�f�>�>��-�Ů���حP������|�G[�� ��t�D����է�aw�} E/��)o�X�н���p�9$�%|��䩃BH&�s�#��D�=\�
�5�6=o����Ha��!H{�m���'T4�6� �.�DJ�qq����(w��N��Ib!�H}���W��[��� ���e �}���[S;�b!`���?{t�PbXFa��w�2䡅~-�52�v�l���������A]�ȳ���6l���� J��yL�90��5B0G˽v��DGGFbOaOb�+d������� D��ֽwd|��n�����`2���e��8�!�����T\N<��BZRxg�q��x>K�)_�z�P��ȼ��΋Ld��S���q�w���� ��~������U7f�Ǆ��X�{��Ndz�*|0���{�S�͕�%��+�`l�_���<ȆF͝��i���?c~?�pgaz׵4�(�ek����p(�jআ�.3��X��z&��Y1�W��^�|�'G�K��u��T�#
��.��7�8�p�hY�r��Ӟ�l��kY���}�19�o��K�F���OKK9$�I�H�ir�F�Q�Bt9����B/pl3;r���P�ذ�i:�sh��,u4Km�W5�f2���	a�ك��6MF���p,�d4�D����b�N �7$��\I��AK	͡s���%�z��@�6R�Y�'\� �ۡ�� ��Nף�F�,S�ᇺ��H%�t�n&6�������� E�~U��k?���lt0Uw��O�A�b؉p��Z��`���� ���|c����H�[/4�g<%-$��Z��۽��� ��J��0q�\�}2��s&Y�J�����9;M�{.�Dw��8)��$���+�peҭx�UXFȕV3�����f���䡝zc��|���RqP0H����X�~o'F��G|��]���nn��jľ,9!A�������o�}�i1�,dc?�B�="�7��\��H�~�#��d�A	���~�J˝�͉7Y�/��98W0�����c_y����~�{�Me�s)F�Nw|�=+��u͉��>��m��(^IN�=��U��D��F07%�V&Z?{,�ަ�"�{�}¡Ё�b��Oh2��p���j�C���m��RwښIz1�D�f��P�OB����ٜ/���s8����P^����l^ZZ����E)O]#x���`%�ñU&�+�o�uL�i�/�&5�VTS�8�D3#�L,�	Y��b@f����w�]��#I���sO�d!�����C���/��ۦ�V������~�l��gŇge�cā�{��tV<Y�V�S�w��w���LsPN#Efi���TN�]ܹL��v��f�kkKU}*mF�0��U��f�7&Ai���B%���yy#�K_��t�Nu����H��KWV�M�����	�ǭ?�$�6��_�et�A(!9���-"���ʟm;�vK��<1;胵c����!_:��
3R�q\a���d\*_�y�����M��s1�p�&��)�y�@�����`��� � }�V�ʒ��+�~,�A	�����/U9?A���n�_�)�v[���#��HB�^�Ë��_`�"��/�������2�8X��)���֑H��|O�:1�qLD��=��*��L�y����#I�&���X�=0o�J��/;R1s�Nns�fݰtc>z{� g�y�ʌ�3if�ʵi����61z�.����RM�rvN�?=��v0�:�
R�򝟨��T�LJЧ�-�a7�Z���LѨ�D4;�U14�bo�r��"���J�ce4Ɉy�P(~Q�a^�5�i�Ŕ�V<�0��ڸE�� �	�j����3�'�]�_���'��ڜYbh�ᬚ�L�lÏ���"�{)===6F�S�-p+49��>Z� �c�"�\���ߐ̜ۥ^���{��H
[þ��,�}�x��Wf\�n�X1�%�jr\�^ ��G�U
�MwG�Ś�e���Zd���t���Y��G�b�*�=��YqZ5qPkOf�v֮������:z#�{�(i�9at�E7Z%������e",�P����(i����V Q=G vo�
7�+1
�~y��U�Q|M#a�=�l�H�b�ᖞb�ɵN������b�^��Z���eO�wn���T]��#�1��%�@m�C��ʄ ��Ő�U`Im�yۣ�wj���=F��`��� W���\�.��/x8��%nt&ʪ�B�}�R���<*+�o�']I�PB�$���o������lH	����%9��.td"'b���I����ӏ�1�6-�{��9�t��`���wU����@\k�����a�ߘ����}�R��j�_�n5�߻m4=����	�
�w*hg���V��+��^��{\��\�G��lI	:�ؒI w�U�@lXf�3i�[LI�����\5�������a�}���M�/�9��R7V�QV	��$s?μۈ����!��lW���G�3�{�7����×��z�����X~��;��!3V�9�e�p����xL&��ʘ��t2&��ovt���L�Oi�2�c�*� 9����D�9ʈ&F����3U����4?pyT4
`*Ԏ>���]^i��a3�躂�������$�i�eؼ��5� 0�����sS�Y��,G����%Q��mLg�����ͽZߒHQ5�`���ȕ,K�����1F�&	V4`$2��k�}b>�c�+(E?'<�w���6�H�C&u �,P.�SheFDTT����  eS���Q�ۉKk�e�-�}���H(���v�8g��s��̲Y)�L1���~�Z?sR��*�����a (��uۓ�'}R�����OV ˞�]N��;o�/�U�7�V$ �"�I	b�1r�o��1Y�A��:0c��n�5*�hy�4���X�V1�⩵��)�iHd�Q�^�I�ߓ���̦p+���#�ޗ��Gs�#i�x�q�Y�N�r��Y�JP�vCj/��S�Kѵ� �v�8��:�x��t*팊Y�NL��mtT����wT�GN����X�o�J*'��B��R�o��_@t�Z�y�Z-��ksy�6+�G�����4ۗg(=P4W �+�W��/���BG��[viX�r	b�伿h�R?�o�T�'�rB6J�-
�@�$�:}1.��;n�)�L��sC��O���c��~��2�zKׁLw���W��ݶS�<�`���6'׊I$�b���Z����	�b�~�X��)-U^��/�xh��� �۔���"Z��=+|Yȹ���-4L^��*9Mm��6��{���W�� R٦��s�1Ȕ�P���y%F���#���R_�{���Wϼ��87#���G2��S�TDl������X|��E0Mt��}j4�n�����1��6��&�ؤ�<�g���D��矷�c�$�$�Y�Ԥ�+��Bt��)����;����cG0��_�'G")�A��%��"&��_�fv�+X}���ab�:[ؠx�D�&C%/g�dmvfr#�7�i���Ubl�*�Ք��Q�63h��O@i���sr� ?`� -��<d�٪:QvI�L1i����X�]���c�;��o��d	)�i����(O$�>n��({�����ғf�@��+G,��ʧb[o^���g/VD� �W��v�=RAW*Wp�C_��I���TU9�Ҫ���۫���;�}TK�m=�,�BSl��E�"1�"�R�	�iVBƭ�-�%��\�G:@2����q�nx�^�cG�b�\�&l��	��8��r�7;(M?�b�E�v������9�07��V1�J���uoPF�bo$Rj���J�k> �O2ި��0��ĝ����S�H��Y�Lt]���z�pmX `��D���$	�O�(	� ��m~�-jέ9��½�w))��?萇���_��h�{@�j�?�wTS[�.�9�=��5
*D@�[(
"(M��H'���(��
H	(H�^Gz�R�B	=���������q��~�x�=����lϜ{g��L�n�٘�@�/��"�O`m1O�f;Ύ���r�u������b��⽨�g����sV�]tH����_��s�
�8�wY�Q3���,�� 'n�� �'�9,Z�A-��I�
¤F-DےS�����1�}u�s��~���^Ǳ�[�����e�=�F�~y4g��[��۳@ً�>2x��Ϥ��Ҋ���7oR�,��]M�	}��Φ �|�FOR� g��U�ünۣ�����qZsk��h�Ѧ�i��X��-���%��W�1g߸��-�/p�����$����}J��8�G�.������gd�(<A���Z��As�d�X*��*`�1���[�.ݞ �B��#%nv�gά�uH�A�+3��P�k�����O'��&_���A��Km��k#�,0K@wR&�[@6�T�M5�`3�UϽ��D�/���J{HB�4�����Q��n
X K�t`^�k��5�@�t��z0&WU� ��*~�z��η��-{�H��vi%�T����A� Kp�t��8`I�:�f,L��%�3��#~z����aР�����7Dɞ��1��5�>��F�L��=�
h�4~{�·�۝�\e��]^$2��\� o��4	�k�Q �""Co\�2_F3���p97�z���*����C����/��*s��6�B� 1��lړm��5�l�0��(�>�Zl�'�韼��4��L����?���7���Z�1hQ��>����V�0(>�GK0�09������XuE)s� Pf�*�]Qq��d��B3�/:b555s@��1ϳn��8�r��3kޖ�b�20;��9N;��zވ����ϓ�+,%V����Ҋz�,�>��L���B u�dd�D�b��V���`���":�\u���M�� ���|e��b�/�]��$,�6j32tӠ����w�whvM7 ��Қ��R�K�� ���~���~��F
Itն������U���X���s�8v&b���A�H�#Yz���{Z�}�Wu�ں��U�����ҧ����)T�@2(w(,=�7��������n�	�����n� ���#p����Z�L򇒌�n�����f��E��@!&y����DZ�~�/�[ �$� �#ޒ\�;��f+'�35�K�K���`�gN�^�7��n�|B�UM o�ǩ�{E֮��a�c8�����\�`���ӹ��G�֓�������Ѝ�������7�
�V�Bu��7*4���p�hOТɫ �Y6��R����
�'�����I^dg��(C��n��~; �q��H04$D����m��
�22������i����p	��nRgg�+���휢���jv�j�k���z�Y���+����v��[�|�C!�
���Pɚ&S�i���nR׎�����Vf�2���9hw�I�m�#�=���Ô3㪐h]
�4����t. ���`�Qf$���#�`��H���Q�[r�T
9��f1�����/˰�V�r5��>��F/j�6�b1��KQ��E�'��,��95yݺ
:��n�&4�E�8��)u@W^>&�V�H�8�/��K��H�O��+ܕ@���)�[ W��k0n�kǗ�Sv~SWW�i	��uie��{=H�XX���:�_�Q�4��mCG��K�3����L24PK�Ȑ��F���kY�"Bc% ?h��.?��$� !''x*�E�x�q��e!p��&X��7���(�1���R�H��h��eZb��&�u�k���������7��US�K^ML���p5�\ݒ�U�>����S9��A�����3���a�~cZR�Ǐ *w��r����[k�m7F�pC���@����^t�W�hT?{a0�Ǧ�K�KTO[u�qp��m"�: |}@R��Ww&��.&�Fy�P2�)h�͍�"\,������#���PE��
���9��[�<�[�3�x8���3�$����j�Z�-|��w�a�k&˷��jU��hU���{h�<��	-�����$E�!�E���9������n�W���cj�"���$�o���`�c���+�'�*�,q�n���ļ�b��ǧ;d��[�)�+��Y��$G��e�r�����}T� Ց�%�ٱ�.�Pӎ�ã<�f�Vn'�Ww���W�f6]��R�4G�[6~҇�s��vôS�p�
���k�O�V�*~�I�����d�����&�#�.	�6ם*�j� ����Ama�H�eR:�R׋����<��F��
�:�?O����P�AË�T���+5c���-J`��+BI�dS�����Z��<^\8Y��٣��TMM��Tm�	�	;�d��Ŝ£��f�b���@�KPQ����$#u�\mӓ�S�<5#*T�U3��S����%	~>R�)�v����"�����e�x�
i����X��H��v�:i~�@��95j���?�f'����V��S�?̩�7�U���RA��&��El��P�{Y?َ�/?��ѭ�v��j?αRe"�2Q�f?e��(��~�A�U*��l���]��Z�VX������� �����RO�z|h���l����O����Y��N�IkG}ۓ��d�t@B�4g��tm*\�u=��O=������*�����z|CP�e����A�R����T�� ����.�kƹV�hΰ�l�,oY������Й9"��W=*@�z���9X�s*���X�)�-df�����'�/8��T]T��|��|�C�!BǏ���h�����<Ԡ>��u�\l���yúQfX�T�VT�\_� �T!C�8�c�n���>":���S1ڭA��g�����h�.#�1�H�n`�1,�g}��E{��DL������9q� ��
�s0�Q�����tY�\`T�a������OoS�Z�+zJr6xxG']���t��g�l{����UH�+L�Z������I�*.�j�V~���
��R{:��~~���#~�0�,/U
�w��-1��Q����^F���⦵�c�Z��û���=�{�6�� I/&M�;r�1���
�9�FU�&a�<;rgbD�`�1
I��}	d5è���I	��$���}� �����[�f"�|���O݈�n>��DvP��((#�1)��G�����.:�'���-X��,�h�b?�$>����:B���h����8���VE�ߡ2�����Px�45�W#�<��¢�e�6�p�PO&�8� ���;�^`��l{�jFur�P+!@����c�d�=�P����Z�3,}��h�:ի�in���Ɲъ�	��?9�JL���wjO��iL1����O8?��vrN:�9T>4�A�v`�{�^�
��%G�^�ގdo}�\��~c$�]�:���k�j:��tY?��-�zδE���i���s�j��UN�$R�U�A�h�^�0��K���[yB�.K�g0R�lfZb����}�۫7Y����+������L^�d�U�)�E>�\�ں�1r�vB�*��HeJR9�
��/� ���P�.�J[�Ti��j����0	����UV>��m?P�|�����5e���������j�(	+;B��� �S�=i�::_
��H%Q�5,6a�	�Q���ѝ���%ahȥ{;ԩ��An�c�����E	����Y�s�Y�%�Ws%�yb��ˏP�㫏W�OX��/ϗZ�焮�-��.52�ϻ�i�'��w{��-���qH]=�k���Po�G�k�l��'�Sb��\����%�& I��"���,��^�nJSY���'��c��DdA�(�,"ɐ��"��^��C7h��zW45}֍9M��Л����IG���'l��d�u�����4��]C�R�Ϣ����� ���A��$���t"�-S;����,g�SJ)�::}�4���S���m�����B6W�4��K�ȷVb���]�T��9� z1!iE�Mܼ�'��1hj�3I��j��?7�.�F���U*%>�X2 |d+	�g^��]O��O��n���s�ǓHǝی��Ʈ�R�uh�g�I	��3.?I���B�V?'���'����&&s��+d;��kx�9��w����e.�='߂�hC���+����ь�M|���)d
h�2�����/u6_詹4xI-�	k�m�s�]�_���֙T��]��g;�xs ��ޣ�����)��$ �̈XC�3V���.K}Olt{'c����\Nu}�%+�n0#f�?��T϶�̮&�6�s����N�n��,c'�/?���j�D�Y�	�ʯS�����Sོ��"W;��C]a��r)���3T�v��Lk#ߓaO�.�4��tk�u5���(Kܲ]��Qû�e,��Q�q	��N���v��nn����d9�D��\X"�v��Gt�~����X+0�>��mѴ}���Qƃ�.�]��8��'����ﱖy~��.�԰m��ڇb��P��W�9Ƭw�^[5u����SexhZ���Y�Rpj���W��Y|�%�\��(���i���.�����O;�c�s4'��߭ �W3����E(k��a#A�	�D��c޻�K�|A��Z���l�U5:�м�����F���]�f��sgk]m�Cx�H�A�M�������\�b�Y7��D/��k�����~%���z�|M���&��ߩ�Pɪ�����mC49VH�2�$P�HX� ?��=cɯ�q;��koT�<�$u���*�8����J=�؍��,p����)M4�5�~��9�h��C�"9;.,�J�:�[n,	Ȫ�%F"DO�?QcrGN������n(�'�{͓h?}%⁪[F2��y�����$a��sI$~�V[�����������[I�y��E��/M& ШR @hUBB���V�U��_�,ñ��Y}[|`#u��lI!�xϤꣾD����ѵ�1N��B߁�`7�*0b�?)��Q�?���V*Ur��o;������&��6�nx�W������~%���q�r�g����}`$�L}��^|������s��E��}�T5؞��䒗��i٣1bAەx}�E�;����c�B��I!��jHMBI	�q�$�p�݉=>�.G��O
|���9�0���wB�� |��IVRn��1q��O���(��GzSS�ߑ��\Y	'��1e��G��T�Y<3�,�E±g�����S�U�.�����VQ��?�>3=����2�O�I�\��27z/�����퇰��	�I����@tl�}�f�<Y(�$��H���C}���М'bߋ�w���p�l��H|=i!��B�O��JlFT��
���!}a��w^v,�
�����adݷJa���uy��_��yw��3��H���׮�Ɨ�,tܥ���������8��ɲ?]�SD�b��O����'����_���O�	���>���K21雔��[�G L})�_�h�C�K7-#FQ�Bydl����ձI��p���X9r�^A!i�>�&l�󱦻ڇ���[�Kuaj ������\Q�Ln�˱�uhU]��RՀ~ f���c�CjK-L$�б��L������Mu����r�y��8O�� ���0���ϭEWpy�Q�V�p�bg�o��/B��,�<��U���z���L>���P%��/<�`a(���ᾅ��L�p�*Oĸ� �ơkR����O���&Y�W���䩀P��ꌹvP�q]�BR���AgJ7����#�4�'����-	;�0ə��)z��9��f���	9��Y3�k�KmZ���jRީZ��.7���gXQ�a����u1R}}b�"�KY�U)>�_�X�u�b�����KI���d��M��uRO�Їf[khXu� ����">�%6�Ay�$���p��`�t4^������+���]kd�n�x�%6���&�?�����UT R<l�jEz��^���x߷��by�j���O$��|���ގ�	���26e��9���rΑA�_RGC�4��۽/h�U�~��E4N��$�À~�/`\���� �W�ǽ��TE~yPƯ�2��]@������W���
�����(��W]���(�����rH�����ĐT��f�����R�=|.Y��e�,�4��O���8�8)t�Ƈ����+Z[4����ꨁ?>�D$>� Ѡ^��Rkvw�q�i;_
������W^��ii	g���O,V�=��R���Nrs?y355�'��א�]^���%��%4i7W��KUX�g�dgn2ִ��x93W�
K��(��LDڟ�<�V��2�Q�
�A4j�-a�����ȗ*F]�0匈�AnJ}Ή�֔h�[���b�9io rF$�U���yRO����Zݛ	����p���mHn�,�~ms_Q�?���5��ncoxwC����4�Js^�>S���E�l��#�d1L���Uk.U䬭�Ʋ�V�Q������D�����ƿ s�	Y�hzY����
�C��;�I�0Ǔ�g��
�ދ�������_lJoj����+��5{zd���}���w�P�u��/���	�X6r��2���wW&��"z��CS��matt�� _zx<%R"L۴�nҟ/��`�K����~]��y�V�H�v��䮏�q���@����=>vQ1�J�b��"$�6���#9�N�*���9)�IP�1O���	0�wrs��/k�cs��;�]��,V�;;Re�Ml| }(o�oh�2� C��k1�c�`���K��wk5�[��^�4>j�][6��8��t:G�io�f�'�C�Ѽm��t�������3�c͡�𕀋����6ѱ:��W9n`k�p��7�HA�6*ʾw���J��4^�[@re1�������)/�U�~6��s�d�^C.X?�S� 'Yu6�{��=���^ޕ ��u�Nz��b�Pᇔ����^�{��9�����Ǿ���������kJX_$�P�����0�^[�f�pQP9�3*ok���0��FZ�N[����]�C��z����9A:�*��t��>�B!ij���x����<�N��ǎ��l>o�1��\t�����6
��?�����
?Œ:�o���[W^����װ��+'��F�%N^�Zu��k���:����P�6�P��=���K9���
^gx�[V\ҟW��^x�Ԛ�%j�;'���C���q��.����1K�*��o�'8����Ú�>�5)>��$�;��ܧ;3<+����V�2�سp.6�I���w��r;*��DL�(����]��2yz�@:�7ɍ"!���u��U7'�t]fbr�=K���!r[䑳˃��w�>�fhA���j+S�Ǒ�
Φ'[����<�Q�(�<Zc/A� ��8=��Jo�y��J�od�W��%z]ɽ8��3*�w�g͝�F;�2�d����-���t̧]�	:4�QΡ���;��R�&�
e�`��4g(�W�{�&�n�(���F+$&[�m�S�|YA*M�=f���U�D{$wN�*Q��O�Jw�+��o�N��6t	��s�N*M]�o��㩶���#���q��▬z�א�ɻ���Ճɘ>Ҳju�.a�v��me,�=��CD�\���kd�8F,�"�LQ���B4}��6�$���qV.yw��p$���T*�S���䗍mA\�{�`��gP�v��P�L��*q1cl�P����yF��-ʊZ+�sn�+����(5���<Q7��_�H+��C�2*>k�R�Vn�%�r�5U�L��W��ԦV=I_��y��|B*���l���"��Ҡ�B���
��J�>狹i���O��TGcG�v�a�on%j����z1fk���@+���Ɖe�@����������>�&����D�^k��x�3�SIPH�n���NU%��BjОd�p��\`�2�`UP.�u���jP{�]S�N!ӂ�\".N!��Y n��V����=���D$Y�>B�}�>�J3��'��/T�]�KP� M�-0��J�$��<?�K����j!��E���ڞ��^ǭ޻������A�5q����i}���^ͬ�F�|c�f�ω'��Z��w"�Y���:3��h�4m�H.)�R39Y��u�T*Te��ګ�P���T5����<�X �̃Z��$JИ�E#�㳫�����	/�x��-W
�KCJ������{�e�a�����n���y�d���<p���z����f�� �:́0������ �}�D��`���F�PԮ��L>��0D8a�\�y<g��e�h�f��?��T�%|�8�2���5�y�_�VtiB�v�r?6ʀÔ�ѿ��d\��jy���ڟ���ȭ�P6�F+�١>��.�ݥ��;V��%��������
��AC[��I�@[����¶Y�ĳ���t���:�����&]��H�T$��9+(�|muD��Df]�V�]�K����P��>d��0�[֗=�|��ZXi�P:�܊0@8�CM5�=�휎<n�A�x"�:=PT����1��ܪ��	/DfI!
UY;�K��yy��5��W�m��1�3ߑ9N���?�(">��LɫUiA���Q]p*�(T׫�S+ז'������(?���w��K� U�h~�e�.N�6�C�9��K�P���T���p�V��k���vC�|�xC-���;��׳th��K���$^�y8-U�YW��L+o�l;��.�ڪ��J ���o4N%�����7@,����q��~��H��G�s���8Q{����ar��ҭ�ϓ
{Ctdܯ�D&{
���#��/k]p����	;�r�7�@' L_T�Os*#	��K����:���4���.��=�Ჲ���J��k����Wx�e3_8���W�;Aז���m7��@�/�%} ��qA
"��	d��_��d ��m�kc��/�yyｯݬ���f{�#4��´����|_��b�Ԅ���썄6q�&��O�T_*<�{:��I�]��]�yk�
o���Q��8�=t璠��S�ow��w��w�n��~\���!��O]�#*��hq-���8�D�C�G�q|�Og6����v�����@�{�;R�x�lŃ�/L�v"d��S�.<�y���g6f�^1���;�E~A�~�%�s!�#U6^��'�˲����U:)M�u��La�fY���k,vU���:n�5�U�����H!����M6�{A�.j���ƫh�g~F��&�k�	؁����)���˽/���b������o�Y�̚����˫hm��������.9دeIn.�F��oьY�r�Q���T���K�3�2�x�-�oJ�O��)�)h(#MCK�+6j�y��O��h�0�뭱T�w~�%�Ծl_�j��8���'���a��U40�!��ܢ��5�����j��EQn^m��Ŏ�bi��`K��CCǥ[��l���)9oCt��L�L�!�v�4kxa�4ܻ����X1�(�YU<����O�
�^�s�C(JkGjX8��d� �[�)�5jiU����ߓ;�_�7�۰1	��(M�76�4mё_$u\Χ�Q�#�&��"�#��_�LY�_	x�������\+�OϿ,����G=�l�բ���@{��+��c�O t�b���涮S� [��K�L�e��|f��{b�q��$�eڀ,���p��n`���`�
�]�
`t�fփfE��!ǋ���7��ц���:t$��~�;�F��-CMSծ��X������ǊuT�_�c^��I�FXu��b}!ڽI����Yk�VFUD�Fl@��Mٰ���k����)�S��6�����>��ᯜe��i�b*�CV�/]��+Jpu�%م.�ڦ��K�Ӊa�7�M1 �L��g &
0��9�-+��S+��Q�&J��㗍����ߧ%�~m��*@�/D�a�z���"�y\�X2�Ok�fQ��7�jB4�[�s�ۚ2��k�r,��t�usJ>�34b^VuLu-�*y�c��W<tyʪ0d8�`�٫��Ĝ�2�;��{z!n��P���c��Ȩ�o}�]{䊚�h $s|`M�R��i+M�����3}���o�%���=�v�M�iŕ\�SV�>?ZL�oY`D-����k9n뙈zG�k�V4���K>ܫ:`�]����5_��=hC��s�Z�Ɣ�y��ŔX�e�Fs�	pV��0�w=�ۥ�@��Y�SE��a�I�&�i!ǜ����n]KXy>\s�ch2�Ϯ�ޡk�1WL.��5�λ����<@�uE�0�Xpۉ����Fv(,P-�@��".\�����\��ܼ��%�<�X1�W*>�C���f�'�n�߽����<P�{ ��[]&
ľ4���A�[y�XP�Lz��XJ�����fu��2�M(ׅ5�A�8J=��n��{-55����[[�����z�J��Jj5�D��+���P�dQ������h�5����"�a-	6+�"�UHTm���Y�y��u�FS����v��<�b9��=v�ѡ=љv&b�q^�I&MZ�0_ւи���XT��e{��5��aA��>� )͸����V��v��go�jD,�� pH1Z�L3�Y׼l�<@Jս.��`z�*�hJ�I�������|��E�I����`�$���w��ڡ��\<��6���}�غ���sA�'$���!=���2o�|	���95��һ!ȕёb�}��Ux!�f�e#J�}`
�O��+��"�z�N���N�θ^cb�)�|�E����Um٨�[B�"���-��))_����f_�3�漄��w�n�c�,�3�vN�x�(�-Ξ�9�"0��e����F���;7��?F�L1� �6����X�YhO K�Z3!�..LK9���g��A���[Q���|��\�#��,w�H����ۿ��ލ����m�1�}y�mÛ$&��q�q�:��8	Hҹ�j���F#T��⥜r���ue_i���8v+�vt��S��8=�U}#Pu�u0^Г��_-�=��*밼�����N�f���Р].\Oy.h ��s�P�h��W�����Eg7O!�}�>
sk��pZ��#ﵬvg�o�����htg�[�G[�|M8j�9��gby��A��������Қ�Fc8t��3/��U�(��/�X�U�5+�R�ǃ6�>�����N��ɫ�斖� �&ే&��4��@�[4���X�-r��+������Bl4c����	�X(�r|kmߴ��pZ�ޣ�zg:h7��\gem���&GGϜ��v��?9HH�n1]�dV�*�o� � @@���+�Wt9�^L[U�KB3�u�Gvyh��-4Ꮚd�T������Լ;[W�fX�(�ƣ���F�k�z5B�TFUFO"j��#�e���-��`����Y�o|]ׇ@��{����ަ�Ym��
cNIM� p�q{�ln����v�85el�RP��$ �<���u�!d�$���HO��44��o���U��+^����Z֟��;;��ywi&[��m�Kx��G��8��ӗ���R�X�9Yd8�����g竑OX%�D�Fɉ�+�.�T%pY�i�;�4�CT�U4�$|������v琔���J'���ͭ�7?�fЭ#U�x/��-Z�X�Xi$�����v��֭�Ĳ�'�"2J2,Hs��hT��|҅FJNMM�:a}��Q���� �[\\�1Z^�d���ǘ`1�! �o����'���y�I�k��j�f(�Ccs����ZG�J{�YE"i�����%B�9Y��0O�]��J�>mh���y�����`O��4��Y#��xs癱���v�C���9Rr��v:s�Wʶz�z8�N�DI��y���snD��+x!kr��&�Jkh>1���tΜ��7ă��E����өa$>���m8��f!n�����t�Rn;��@���iGb�9K�ݡ�Ϳ�%��l5l�mN
�+/^�F��rZ������4�#��}E'� ��\��&S'��n�y��lN��Z=?�����cY��X��� �IAN=	EW)�G %�BkP����P0�ۤ�u������'@�+�v�lg��*c��F{h�p�{��u/_r�a<ދ)'�X@�I�����U�����]�n�2򜎔�+{W({�N,�Dj����O���B�����H�qJ�4耓�:<@S���f����/^\���Hx �e��ܱ�'-��Íh��H�M����[Z�F�2�۾`�]f.8��m&�ݭO�i�̖>���ѓ��ޝ5�͚ͅ��ꐎ�]��A�ɓ��-�8�=;;�?������*(�/9`@�<]�Y>bٻ����=Z��� 	S�TU���!�:Kĩ�����9`�ڻ���@�oO�VK��v� ٹT�r��g���0��|�j�~v� ��a;��\���.y�,���6��?�`��:__	u�5c�D�G�}���Yt��T�$VC�r�'�F�l螬�[�nS�B)� :�!#%�+��e����� 1�.~��=-�6)z�Mk� 'X�Te=;@�a����	���˫k�x􆕫�{�n�~9����G}��<�6$,�f�	WZ[%��׹��\�^c�z�|�)��S�����x�Hm�����[$]z���Bl��p�R9��x_�sV�Ӥ��i|�]�щ�OZm�[����U�Zz�Ǐ�)�������n�*j�� ����m�R�����66�ݼ���S���Y�s1׳o�QF�s݇6����y{+����)D���s�/+P� �N������K��:^O�A}P���ꀏ�ޯ����޼�]���F��etg����GG�u_u�Qd^YY�zIC���g��� g����.l]�Fo����#����hWӸ��ǝ�;�$��?�S�\O�yVn8Ja2>PefͰ�\e)9�(˸��8�D���j�azz�
�E�-4�Jtn��Q��]��G�"g��$�?�@�s̺���?����/�xu���:8��S���|(ݥ"_�m�qR���	͸���
M��:,�v��3�QA�|���P�4�\4A�h�{�w�;�;j�]�47��.��X�e5�40NْS��U*����΄꥗q//a�XB�lx�X>�O%���|g�@��Y�\��=�{"fD��G�΀bM+�%���W�dS�ʕ�8z-��9Փm
��.mkm�~<��0�1]z�Fd��_��~s�*�#���B'����~��\::���I(W�+X@R
�jWjOAA_�RE�'5�w�*q����Țz���]�%����1M����7��[��s�[>����k�{:2ǄsH;J���"JmO�(W�'O����TSR�HsDڕ6'Q�Hך�Y�5�l.j��$����<:򮾈Nm_������O��T����0�0B:�$��[�E0���r�$�mz�pIIiR&����M���iڙ�~��W?����/ƆC���S����H��%-�)%+�
��K��U�is��ϊZ�X��q۹��&ݬCCC��w��ĳ��?wa��W�{��Z'�1����y��THGW#]��vM$�����6�Ji����
e���T��a(X���E�(�n:0��{P�����+"��g�6���@W�IU8ûg�1ѷ9:e�cf΢+�K�'�6�%"]��띢Lq������Z�H�EHx�؂�u��՛$;}թ���\A�S[>Y�[X��6����' K�t����W����Pz�P�.��T@��������+�,�R����ޑ�\�=׉=3Y�M�w%V�~�gs��Sj��O�Н��W�������X
z}�DA�V��"Q��g9�� �OǦ��s�ͣ��#>�֒���í�'b����{�}/����E�`bo>:|B���ρ�/�k�կ-.oV���SQ�ÿK�K���P�n)�It�P���ĺo<}�)IW�V;$h5m�����z)3��>�۩���C��8��s+XI�5cB�W�*U��/l������ze����k[��Eih�;n�vj���ߕ;Gm�$���-���u>���������s�~��y����p����� �8T"��!���7��?[���}��/�`��g;�9��-���Ō�|��k[;}C���O6�,\��iYJc���x-��j��������龧��U���
u��z.�8���'��p����%˜��`�{��K��-Z�y��ȇ�UznMY^G�&�yl���E�R��X�4���w�·��Α�`�A��8��fjE
t�.�}n��xFz4�������L�NE+��$�W��IC������\�j4>	�e��y�ݬԽ|�`-��1�s�d<������v1A��k��~����xJc�uYɃ�Ur"���%.8��@���90�g�D6]�*"8*Qhl#�����Xln���m�Xf�֩n�k��&���{N���ͫ3+��k&f��>B�&&E+�Sʓ�$�0�$&��(���ǯ����L
SfR�*���H��ERP3+���K�0ԇ^C�� �1'��K�#�MMM�3s���D�&=�i����?�^ЗyB���	�-*2��^]u��}���_��6c)�x���
_oŊ�T����&��X�����Sv�;|�?��W?��ϙ���_���_\��W׽�	IY�MbFb�����{�hZ��Ueܶe=��:G�C�z�d	[�Vcs�,Y;��l9?$
*�?��o�ϗ�����S�[�u�`+׹�\P�ӑ�N���b6�er_a;��#�ݺ�r��5����~��G�D��UV��6�~}��b�
n^e_%멃��4�^��z����Q���E�9� ˮ׆�Q�Ha�Q�K���:g�d���du�/e�׃\�/���[�M�C�V����;����ʾ�eԚmj��%�?Q)J��h�#��O����EM/�(%�J<��[e�ᢰ�֞�׾�*Ŕ�����d��-��?�P�f�i�6j���?�L��ea�fev{}�=������n�3R���y�[���n��kf{O���}3��;3">*D=ݶha<���_��>��9�
�l+((HZ�g�Z��j��>�m�%h�p�6Q��c}y�l׺�5AF�o,�B���#_�yv~�~H���?����vw�:F}�J�@��I��9�^���〇���$����r�٥�s�Qc�%��I����!;'~W0��UDe���ͽĆ��ӓ�QV��
�d#<�'�y3MJ�^�R���t��������}9J94�~�t��#��.��C$�3������g��nf��R�R�G��u�r��9f�F(Ok~.?�!�[oůlp~�������x|C�����Y��.�����=�uO�	������P������'�&�⻬m̈�sQJ�t���ݹ�I;}v?���?��?"�#���H�)zg���ݾpH��jS�1K ��V�P��=Hw�l6�O]1J��He��Z=2���tj���{κ�ǟ��7�v+ܔ-�BW[?��+'I���X��'�׼��>��9f��:�m�Aw|�x2�d.�`V��ĥA�យ�(�@_�%���.��,"�'�o�s�I�;0�[���1�y>�6oQ�U%���.���[�C�t�C�=�[dm��E)��-��#�*{�֖|(�L救�xUS����$�_�P8���[�;���iѩ˧'�Ӷ*ػPiB���'�-�|;�C���-�2��t�`prk��1��@�I�>�C�a~����k}�)om����v����Ob�P��דs�`\MIXw9w��6���#�K����&==�[s@w�,�U�9n0$�V\Μs�ۓ�{�b@1�[��?R�c����*u�OJ꘿��6+�El��۬�=@*W���҈����O����DY��y�Ċ��ʷ�����x�Ͱ{s����F*b�n]�����PtVn�+�9�����Ğ��S��rW���}~E�_�$+Vl{X�\w㪼�����xM��0"Xtu�b'�����z�uM��z��#V�>B��&�:)���ZZ��/<����D,�Dqf�ZJƅ���)��6C*�x�gVz�����Yԛ[������}�oH���=�A�G[/��8u�/�ۓ��ƶ�+������ ��]�|g�*y/�_K'`:�WfV����׉�a��P㇎����e�o����Q�S�R��(�

{����t��-iZny<R|�����Eov&�I�������.M<��6�n"
(i��?���9�����"G�}�[=e�8�Bt1ia�ma8�ͅ��\�F�_�v�z���ˇ�_:n#�O��S��s���Bh�[R��?m��:��o�?NH9!��Meke�ez�2�+6ce&��bg�3⳽��+�Ҍ��R�k�$/���~97��J�����߸�Е�s��L�������MGRz���~���vP�v����������)2A$�ӑ�n�ª����N5����r�����o{׸2�AŻ�I���tmy�O{�<�m-nxm*�#�,%�VUs�u1�_����>��U�V,:��=��ȱ��q,���_2<�"�V��#���#m.d3�:��Y^馻,tt�S�itt��=JV)�r�u��(=5�r>���C#L-����&߭�?�m��KܹKmh'�6,�sN�H����ҝ�m����{\T�Ua���������Gz)��u�D�
�?zq��Um#���N�kV>�g�Pm{%������%ir���b���f���C�|��J���׹�+U�m�v�6�Y�K���N�n%R�+�K��JS���Q����R�Dr,8�'ń�0��e��D�bj�*+	�&��2�������&x/�jdk����ֻU1��7ݼf6�[!�m���z]����C�����_#?��F���Iz�P�ܩ�j��C8vc���-o�EX�EU2}\6cd#"�w�%|�N�ן�������w�W��bB���޽?�;� �N�h��UYZ��������EM� ���թ�����_���AOؔQ���gO�~�wArT���MV,ݫ�W���,��(����<v�O�ɑ/K�w��)����I��E�t'��d4�"u��Q�1(�[hq��/6�ƴ��|���cbC�犍��8{_M�eդnz�L�A�a��� oL�K�.���Zn!��d3�_�(�0������_p�i0��;iӚ�!R�l�6j�༉�uH����ߗ�.���e9���u�%Ň[rž|S���%��~1Օ��{s���kf��sk��P�0aD���2_���/O�}�cYW7�z���J�(���e��K�ߑW���c7>n8��>��;}�|�G�]���;��.�[��O�������?��
�E'I�$9v)G�.��f�k�<u� �[Ju���q������Ys�VT�[H�Sf�to��i�P��/�9'Y��K��Ysi2�r���ٔ�]=rcX�.�9�)�\�L3BL��?��;���}���bAQ�bDE�"$4E�w�
� %��F���HPZ��!�"EP�z�PB�3W ��;��s�8����1₵�|��>�\s��|{f1��xx�3�|��x���3|O�iG�B�8�m���r�'�H�PG�ʱ۞�.I��Q��W�?�[+�&�Rb�`��+%�rK�x��}�_��.)ﯖ�A�9tj�̂肏�F㵂��y����1�4���O�,�J/.b�H�btuS\�\r�aolұ�q�艜�������`0U�T]R����R��N`�!���	�g�	i��jfƹHV_�6:�]~��z�3�2�g��GI nqR�#�Qg�2��C�2c�b���u
�eA
'��U4���eϸ-'|����E��+������?��/�k�?�D*c��[����ѥ���c�u=�Y���R���C�t� ��4���7$Q��J]Ӏ�6��)&a?]�d��`e�%/��.g�5fae�Dc,G+��~!A�2	-I�����r��������hJCʺYp����C��o�S��U�I�A�J C�E�^��/¨p�˅�.��u`��**P ?"z�/-2s!�y_���qE���ɶ��aݜoB��:bhQO֍�ṷ�A)�S��"����,�E4��;5�;Yr{�������dN$r��<� �%���K�i���N6d��w�}��x;�޹v�J)�Oo��q���h���~e4�P3��� 1�;PhL���F�j7�$Иk�loT�h(&�Ԥ���}O�g�ꨪ+��} ؑ���I��Q&��Oe犥���bG�mV���w4R���]꩞H��p,~;���q9����O]3^����R6���i@��<r�y��,�RW�
����:������G�{�vkn@�}8���*d�G��%t�[M4���0���xO{��<�IYf���#RE��u)�O�2��Q��o4�尿�%6�#�֭���>HJ�����
I/m����s�ט�s�1ӑ�|"D�U�˺
��(n�TF�7]��`���N�z�7i(���Sq�ֵs���X��҃���׿���{�K��K//,g�:j�1y` h��/��r4K�r�PM���m4~Fc�GISQF�㸨kB:�}�;�/@)ʛ��&fd��0����e�
�**ǷL��{+���x��8�h,,sA�=Sc;i�����#�&����J�W����#��U��0���n�y��V���N��w`x��6&��p#�i��z��<����*oi�o���_�w�_4A=������>"�^{��/vG���/���b_!����M`����+a�]��_Oz_��y��"�]�Sxy��G�������'"�Ul~3:!��+0rCc��R�N�7�r�/�T�r�&���T�괛�~��0����C�J�h�oZ�l��w�,��/���2χ�p�ع]��E��^��jcS��jR[ӄ�9�lK 6��.GT�l����v�1�N���R�g��չ̸��	 �_t�U�����,�7��Td�{�zg�#y�0���S��7�_���o�8�
���� �h�W����<弴�Y�R4kP�h����@f	D��=IIzq�ɋ#�_�P����6��2��
���W]����_��7�t�C�7�u��+�h����;�N�dN��?����@���F䩈Aޱ/���������|�f�ς��l��3B��~�ȋ!(�v�<[�D�n���AvW�/{��V�W����@C�<��y:C�3Q�2
�Q�"�So���=Gt�ܗ��2B���Z.��� T}����B����&�<��V��";��?c�4� �bW�]Ruv��Ի)��������ޓZ���IR�h"��g��^��?P���Q�ʗ�O����o�� 1���"R�_d����q�S�i�uɢ�{������N~�}�"�Z�X��W��u�Cc����{��-C��9�2ۍ�OǈK�e��}��\ 
�l�'/*ۊ�ك��w���&(G��[H�u�t���Ŧy�{�L�by��,���b��x�\�jSE*u�Rn��
��xI1������}"쾖@�U"r����A�=R0D�X��M/�$R���ݳ+ٓ 8�d[��d[j�}����#��T��^`ey�1(&!����9��2�H>Ewz��X�-M�tK����Oɇ����d��LN_p�Zv���v�nn!��ñ���^	��J �@a��Δj/�Z�V��j��8�~.]?���:�V$���)�Y3�l�a@Nk��$�r�z�a |Dws��zv��r�cs�g�
��oQ��J!3���K��+g���Q�]���oZ�[{�� ����{���M�s��|��\'~�݄v��'�Jy(����Uc��e���i����_db��B!�;sW�{�v���x����5�aU��2�}�&������Pz˩��� ����۾*oh�]{p�co��z?
�;��IC=�	��	������ {����Z7
�Fr��뤘'Lh	����fC .c�DQB�Tcm�'����'N[�LD%&���
SĔo{��k��>�9=�0u��JWJ�eI��=��z}@����Hr��Ձ
5��8��c����4�c�/,J5�A	wk�����Gd��9���� 
�Ի/�%�@q����2t��=�󏦅����f�8��Hl�&��n��.OWX���s]UV��^���9�z�z��~�F%����IK�}�d��	�P	es��/��L��d�We)\5�z�v�ґ��´�c�A��� k���<���~�W�����Ꙏ�f4�9�1]�$}��c���p�ƲT��I��|B�k�YM}�༃"r��ɀҁ�a}�""wc�7H�p�KzQV���9z?��(��joi�΍�sW�f�%,�N����j��O�I��O��������)M?D'��y�c'�ͩ�s*\ Ƹ���>�'?�t���2��H�G�$c� ()p~�N��V��`nc�R'�3��D��$��k�P��^���&&�EJ%��CH5�%�V��ӡ�E��c1Ά�٠���2=���%ÅrdJ�����3���)t\��C�Q���8 ���a�,� X~��^�@v=�
�����f���I{�}��D���o�L�\��P�#f}����9-�EG�c>����� 9ʋD�E׹�nD��3�c׻�
P��j�~�X_��sP�*��!��YU&25aL��r�eD"���~�U���鹯S3�p<���P-w� ���~�������(��Oɇ�k��U��:��C�~%�L�0������2�������N]��<�i-�9��;ya��94%]�.2 ���D���P��r�Ʊ�etN�S��q�Zɮ?�Ez6�����9�
����6��b�'2�_��������+kH���|�5!k��hV�xƧ(Ue����S9��MO�Q2wUYbV�T�2�k[�[���R�90�Ѡ0��P�~-�v�&c?�ߐ:U1<�-�8��*��$W2*ZΌ��9�
��.�k�������w��Y��M& #D�¥,��q_�^e���2c�s?\��4�?`��\$x+h��Ty��/��6�I�"��Y�5w��D]�8И���}���l��Z����}+���Uf9v%�����2ФQ��̔�0��t�:TT�,���h)[������=�y��c�� v�����QM{~�h�KLKoG�P����*ui��T��lU����ʎ'z�]�0��0J��B����Ť����ZǤ(DJy���a���)��RoM�o�w��(gP�U�6W�5bC�ث�XȰY�m��</�ܷ�:�O�z�NS���ې�Y�g�B�QPR-lK�Bi��Z'��z�=�r�3V6���V]���\Ա�C�y��!�fI���kH��>j��o�u�#�4az-	���p)�\�ei����V�5��O'����eȞ�Ъ�������.��	��������d=Lο�x��2��i��/�����	*.�������IJ�\�K	�bD��N(��N_֡��U��!+%=�f�k �m炱����B�0hԠ��Y#,{�]��4�0\ )wx�������^�Ѓ�fZrHx�*S�e�kŞ䰃,�Z�P�s1!mǷ��g�Hر��1�����PL�޺LN��R+A�R�a�� ����s��`��g�����z2���"�-�afy�bh��,�o�h�YZ��b.��]��{����x�1��k��0�3;@�n��FOf到� ��v���W�86jy�I-;�3����~����g8��������8k����+��_9��_�=���Y��|�H5��=;�n�SX�����dGt����i5�@8�Ж�ިX���g}�캈��h�R|����E��J/� y=V���aĮܵ���x�=���y:4?�T��O�����kǎ�[x��Ž1���pw_:�q6	�迓���#��]��ݗf��&��IE����^���B�aMK0D�#K���2�1�k0�ٔ�A_U4sb�U��*6��M%BW����Y�4N�.�	���m�_�b+��q_Ķ\pq|�N�Ǿ菮��z�T�.�	������ݴ&�UO��k�=�_�AEu꿪x��%�P�,s���$�p�y�E��V�0�oe�b�oPm	��v��?Έ��V����^e���:�������%��5���8sC\@�L�\�t·\v�1�|j���>ij)�`>W+���`�k�D��-S\%����M��eC�)���c�x��%���Fn���R,'���a��-�`v�#�3}��3Z\�Gk�e1�a�l����gT����>���q��n�x�

	1��{�3�{�]��9{K��	�@��
���M��O�/L���M���ύl�.E�bS�� �H���9jQKDJ�ne�U_NX�}��2����cc�����r�r1b	X^^.~2��>T���=��ʵ�\����L�ݯo�-T�DˊM��ފ�^i��&���\�Da�'A�$K2u���mֶJ��-12&&��1�7���/e`��?�>�S�e�Q�Y�U�V��%8�_z�1�����U�|T���ux7,���������j�F�WB����E�����OK�������?��?��������g�حm����g2+��8���#(�+1-�H��8>B�B�UB��2�hהPB��3����19�E�;����}E�7>yO�R;w/]�'���K��h���>�\}�v����/ND���(�r�4��R��r�N$C���T �m,|��v���R4L���фM�:�>~�����7ω�4�q��n(.�֣[���պz}���Ob��w�-g٤�c�����Xf��q��J�i������=�!�����tg�;�����A��c�l��y`�]e�R/:`\k"YT�|hX�/B̈́4�����jω���Z���m���&�ض�����[Ô��ݯ���z����ve*�'�w�^,����N,�~�{���AW~���� ������OĖܓ;Q��ЉC�.3�/�+�lj��1�ؖ2<����A%�/����Z�~A|e8�D��LWqZ-�y+���Q��/�1����Au�:_9�3�!9{�b�d����婱�@�lG��n�
��7;r;���Z�IԾGl,3�H��?�!���O�C��Y��Í�oO0hL5m��~T혐�|�5�nT��q�[�����YY��l����O��}�6���t@��O�Z���P o�����g����gr��i��ӟ�n�?���D_/ ���D���zg�Z�idzD�/�u&�/�:?��Ոsē�����hr�,q���y�c���αo�ln����fb�����;�����XqJ�L��?��`4�_�@%�_��������m?�%�
*^
lGh��[�T/��}�_-t-|��x��2ڸ(��Mb���r�����OxiA��s��M�:�G	��ߓ�
:���mL�IO�{�I�?H��tR��
�6Z�G�s�	�Lm2#aY`s^��C�6�i�Gy;����U|��γ��Y$K�����6�j�=��Or~�/�����S���%s�hFOX����c���x� U�����?��g��I1�4g,;�K��#��05�՜)�To�"B{Y��Gzs3j�ú�?��[�6�u�]�Y�9����Ũ�a?���me�]]��94�9܅F-�B_��h\_����G東/_'�i�[�x�)�rn�Mͻ�r�X�2�4�q��%�/�f�y�jH�"�Mz�
J���l������lR��_�=6�茺5i&g�LB*uCg��0�&D�hY�S��l}��VA@��D����>�ͥ@���T~s�}��މ�tx���p���q�!�R�٩7Ʉ��J�7���n�Ն��S�~��8��aR������m֬�b�~&E�����rq�g�C���}u�W�j&j�O�;��D������zr��o��H�(�|������il�;�-��}��w�D�i�X��,���W��mwB�ܜ1�9e��[�^�h��蟏$�k&
g��YD��X�"��q���18�z�@,��▓4�E���܉K��uV�T���N;-f��f��oC��IO��[>�+�a�t����U��iA�D�[E[��jh��ƣ�ԋ,/w�寐BZ����GJ�5z[��>�TR�r�i�U�>6�1E��ǳ��(���כd�:�)'a�J�V��s��jN!	��:{!h`k�x�$
��"U�m�ơh.[V��X����ΚM
:f v�����rS��6���w�-ھ�/[�/jJ.1�GJw6L�R�RUWf�T���6�����X��u��<�����T�9����XB�2�Gٙ��؅Q�U��
$� ��7����@ qY�l��/o%�D�P����X~�Dw��h��w}"(�q�\ջ+n��-HǋhLfxv $?��Й���D����1��Fev���.L̀��A�,�!�����=>,b��AO�Z:c��}�M�^��1+�U�ՙ[�RE��g��ތ�~vS��[��T���7J��l��.���fqȷ�2-*�iRC�{�i�1�������8��<��Д+_�v�E'!�A,���e���ȎL`�J�\���5f�¯����/t1�?�R_+��+"�2�7�s`�ki��}u�.��.��K�b>+e|���&}[�h����V@�א�p՜�	����.x��z����i��&_��\�n =��.Q¯�1�OCe6�}6]l�A����ͨ<�d��1�p���bS��u��	;�kS����������������W�1���mX#'�`�r,����Q!Ĉ	{�W��Ȱ��.�)�$ljz�˗��y��S��l���1{(a|╰f��w����ܛ�3�p���~l(�rK��)��N�l�mձ�K������R�h�3�`��a�����U�rub��0�!�O�+%��}�̊.ݠ��B��[�(�F��(Lz/�n��T��2'���Phk��$ ˽����!�n�ܯ5"Ν�fLpXq$º͙�ax��v��ծ�~�|�V�9òc��'?(��
ԭ̱�*�8N���6l)�=9�B�0>=9�3H�V�R?�z�%�K5s$7΃�I�B�fj���V�N=���L,raAӼ�
�x�a#S��
����q�Hi��Չ���߀p�Kq��#?��vm��LX]���=ej��bi�l�N8l�ϕ}�q|8&|[�?H�Ŧ�G�N=#�A�Y,�OK�u�x��ᤸa*���?�"�mH<�m�s$�)��9�ߑE7�����B�Y��S>��?ĝn�-��A|�O��r�>!�dN�L��?�^�<�t�#m�G~(\�+�E�x<�~.�<{Ǳ)��K��O :?T"}D���p�\��y�q�T�o���ʛ�ג����shu�W�'U�s������5K��<h�}[sL¸T���hB�Z(���N�D��Q���T�N
hξs��s���/��;�&��^�}�Z�a���3̨�o��=�L�
�{ç�*���۱Ŗ<�u�����%�MTM�Z=�g�4�!W�P�)S"z��H�{^ϓg���1,ŚI��'ɩeia���nB�v�-_�<��T;* �}�#�M���͒ח�}�?�Iռn& ��>����4P.4��h��@I�![w��9���^�`��_CD�uޖ�~��70� ��!&�2���k��}!�~�I>C��᛫��gyv�D��I�q����m���[y�ՒϮ.f��5ka9�,%��t���x��(0��C�*+",��=����0CW� "Ӫ��ݮ�����Ge�Y���q|��g�A=\v6݋���N��<cm�RۺN�ٳ��)C�pͺAݞ ���[�V���S��N�!�~����e��_�a����>���z`�WW�+
d�C��!���~����%��� f�VG�(�Wˤ$�/
O�2.f���V��W��}�k�Eԏ���UgD:n@��a��~:���6h�ϯk�GuZ╎��t5�T,Tcy��������Q���m����=k��4��9q�*3�_H��q��c;��٦��,m����(�
�|,s���e�
����2��X8�0H��Ɉ�KHƦd ��jvSVU�G~���CZ��eXE���@U�{ٔԫdP��<��~}
��k�V�釟����d�3�|{��{
��?��x��ti�o�l9��3{����̏���R��vp�,�Cy��#�\��{���6�e&ˇN}�ed�춭t��.��u�6�K�N�4 ^�*fTw���U��u�詚��)�*���<�s�����F5Mҵ�܈ j�-;�h��~	�OR۔T�)'������Q�khL����"#7M�u���Hi�ڹ'c��=+:?��z����U��Po����.)��ʵ3�<�<j;=%�Z���+�P8hFup˼<o*1��$�q�*plUPFZf4M���j�,q ��26�b�+�@�a��[~ئ�c�m�U�R_?tt������c��!LB��9h�D��je.�!����%���-����M�����{��t\��V3�j�S#{�'�v�5G�<�> ��u�%=K'N@�o��^�_��&�9�>҅R���x���B�js�04���O��@qҫ��Ɠ���J����7��Ep����	��HY�\�j��Wq�^��_�����|�ٜEZGvu�^�yڻ=���4���Z��[Ъ�w������D�� e᱊�=%N~)���zji,(�~�N�t.4�G��M4����|�\8�$�VR*�f$9LX���:�4�0���Dn���R~���B{_��̰�� 8Pc������:fͣtU��NUULps��(�|��w�`��[|�!%���~��aA�p
���΋nE��[l t�cU��׹�;��ih+�y�@�����N��[~qPϥeY≰��
�8�Yc�$&�؜�9�kj�2�K�O�SP?���T��C��'P;�sD�1G�n�QiIr+�cU.�B.,'���uU����nb�\\Z*r�� �Oi���
h��0[���Pă���WI)����F�4`�n���L��Oƿ}�t#!ͧц��}l!����Ufc����^m_��Q�����@���� D[�N����#A4M�-RO�Y��7`yO��D��(���6�-�F���HbR��|b����
��+��g �,K��:8p}����7?��0��]˩MGa&cu��Ft(�j�䇞������qL�ӝ�t�ya���d��V�`lh����Vg/=�́��$(���= ���2X�k�o�)P6��ޠ�7i�-�+>�ϧ��a��o�.�����Y�i�����R�U�Olŵ�N@�kG���0Az�^(����XE���?��zS~+v*�j()&e�(�A�����nn!�>��j*)0#�s������a7�x� ������̉����[��eC�I�xq�T-SIY�崩c������;fR����sm>۔H_zo��_`u@_D������Ƣyކ6�QfH��޸��TS��|#띺ܹjt[~�o�Y�R
�Nu
a�Tj�� ����K.q�w�&��粼(��p�N��O'� ��Le�'˾ڔ���eϦe[��������#ݓ��Y�t�UieP�t~�'_�B�B�S������	x}z��)�U�8i�Nd(h΀
1������sQ3U/��"ʽ�L^�d�7�K��(����˄���&#�� 7��m�g=ס6��^*����`>��
��V�9�̷���&/ٿ�![��[��w�!:	���t��ƚi5I\4�E�9����d�n���$�'�ʗ:Y�bퟺ1�l��5�y��ħl���˻4�JW!UNZm�mu�?�� �(�JV�Rp8�#'\
��,�6��Hf�SF���x��]Cg�����R��*hIjK�Z�̰N�W�@�I�z̷�H�b�⍟�V	+Q�-�e/��U��g�������;�H'��e^ӱa� �i uK�_�~�B�H�y4��{�y��� ?�q./�u�_[e#�R�#`:�E�|�a+�~^�R�@4���� �D�=:�WPc�Ҕ���ضP�y�TA��n�h�S���a�qu�t˝�*m7��N�\:䷥d���+J�C�Pa�*\I:tM��.9�y��r��ko��	iG�^�7�w�N"�ԏ����}f��j�Y,4Pz�3`��A/��m�
����ގ�� ubL摫OK�q�dq�J�CT�/$玲����Mb�g���
͡�YR��/���/mTd`7�n��d��xP�)Q�W���ؐ�wo�����9ض�\ ���wS�:Xji%ᤲ�X��-C��wÌ�:�e��U(߁����%�?��#�y�iׅB�� G�Β��|�`��T�TGR2�{��j�-���`�h����:��ȧ�.���C������P�˗�׍���}�~��xt|l�Y�9���c�!L�cIs�Ҳ0�;�[��2���4��������gQ�����s��1G���D��>MR��۱9LS��`����f�|���	�Lʓ�UG;��;@�q^�4����w�|��+I�.�Ѧ`'�ZͰ�g���$@,PXn#�-��蠖H��	b�:�[H�}��^���pQ6��������G9�w�*�`{3yh��^+�8)����l�.����/�a)\�]�*�1���'��h�i�A�SM�X� �vt�@�%�k)fa�Fux�kt"1?1�u��pV��Η'���Ql{�Vڷ6^�&�B�[����g����+�F��}w'���	e��*�~ЌY�5������z�Wf1�uy�E��s���?��6���XB:���  �uA+���7�����+G�T��a�J�+69��y���!*�ѽ���I�J�Of�a(�\"�͡�&q��F�p��>}�jf�H���|�18U��DfbOl���1�(A�H�����V69�G�����k9���?�mh3����~�� �R�zM��	� x�k ����@����GuѺO�D2t��m�8k�t��mщT�Ԏ,�p����5ӎ�<�mX�ba��6tT`��J$r�v7M�(��m����"�:�����u�a�2��{�tSt�|"6����EM���9�-s�3��lE�+����P�],��=��@�%��e0Q:�~gށVtr�i_�IKmQ�̪�C���OȌ6"o������X�uF�zeB\N��G�D#�c�V�|�S�C��m�'��P�'���7��u�C�2T]�)�~yX�R��ab�x#A�Y�؄�����Ne���Z�.����8��?М~�m�8�?���:�їc\�r���\V
�إ��	�5�^���m\v÷#4�_	�Eԍ5	�Z`i9�G�Q�I����t�o��d\�i�
k�C�����b��M�iuI7@���8?�*g)�<u�����6�p��G���<=�� 4xg�ywM5��%7��4ԋ�1�(���)tnO%8�d���d�l`<�d�4��!�;"-e^bh�:W�s��۔3�h�e.�L���������!��LN�*u_r�oR#����z�9  �(��r����<���Dv"��)k���~ꑺ6����PE;�Qr����q��L!�ۏ���Ay���H��A_�)��&�l��w����I�M'���PQ��f��\�XN@o[��<�
��.����"JіD����bX��:�`}�n�+����.wծ����"I��m�0��®pZ`�u'�8ծ�i%1�+�[�'�@-C�Z�����e<�T8�1E����X�����]��u�4�P"�!M��k�����{�n�]f�	��ֱn��ׯ�Y��"�*�>���6Ƈ��D >x:�tbLї&����A�8>���gh��vf$�j�����itYQ�ϙC꼶�F?�zkZu�r��Nӳak��k��,����d����v�h�"���{u��bϽ��������Q���!�����Yi�)����~�l(�ӛP�[�"��[lr�Cy/�F�+ؤ��6�sJ���;vN�Ilz�ne����U����[�	�[V��)��#�ޛ�ei}NQ���B���\"m}zNw���`�Ƥˢ��ո����>{w�/�� �,�J��]����C6vLUp�p��A�z��ą����^[T]F���ͣ�S�M7J+��T
+3������p���u�t[	���|agjG�|Lh��{С��xoa]��"�J�Do������;9�<۽]󳶞�Kȡ;;���.��z�ۄm������UO�DR���[_p��\��Z��љ�3c�*S>�XyjtU�É�Z!��|sɃЯ��<�1#����L%�Q���Ȧ�iR<�@n��uwJ���V��t7�dt}�v'�(u���3���;ەߘ���LUn1宧�����26����W��Q��"�s2���x�׈�	qƽ���e\������7������l���;}T���,L�_���ᰲՊv�<���u��u���JHZ���S�Q������."�]�FK}Ɯ���P�C�%��35�V��#�(Ƕ�ve��ں����%j�T��o�������\�C���$Of���=�2Bݠ���PO#)�z8i���D������X��Z�&$c�������V�����6�,옍�0��U
8�57ֳ��?��N�� +�-��	��4��R��l����`�/(�mU��6/"	d~�ݾ%��rw�왱6@ҫ���L-���B�͔�jM�F��ׄ�˼�ݎ�'��]{IR�5�xam�Ys�4���͢j���3H2� S�6���p��[n�J�B���sl{`�6�9r�J�-11��EҚ/\\q�1�u���C?{��pS
�xr��7_-����dn.	Ҙ���U�8/�:�l'��d��U�Fw�er��J���?��يl��P&}b	��YX%i���fz�,�������.������Y3�sU�%�>�j7��Hh5W~'6�)��Kuh
�N&�����{/M������C�2�"����PE#��=i(����b�d��W�Z��/kG���
�9+9�a���H/�����*Z@d�즐�v╽�PDy��/�a��5s���m7(&)�!SAz��wy/_����{g�=�	\X��e5�xA~�Qw�S�����O��p��`�����B#oV�V��R-����(3�읜��EE�{+�z��Ā|��k]WT.��ӧ��k,ct@b~���g�WPA���m��/ވ�����Z�T����mb�h�lx��3�:��*v���6"�s&
�bǆ�C��Y����f��}��F(�v��v���{����,�������|�SKcoίz_o"G>I���5��хNc�Cw��0	�bAm՟_�����$h�[Fr��{�MB�i�oVlͷ#,p��w#�h,���<c���H���x��M�}���]~�z~�e��>�@��;�>&3�k�u��T*f�bt�^�#�xv��b����bE~z<�O�©e��"���Y[oM�F~��˸�j2VY��N�bMx��l�Wmkh�Dm���p���� ��!��{a4僥}� g��Pg��j��)^�b32�a��w�t��M�03q',HLL	H�\[b:�h(��zR\���;}LS1�b�Cp�U��\Ut�bݤ�B��EU��:͖�kQ������5�e
����?`���S����8(�<BV����C���ǝ�z�d�5���&_��	�t|4�łH���f�Ά&^��k���U"~� Շ���X�ʅc��i���Z���i��Z�R�\�f�g�]�>��O�~0hEsg�ě\ߦ��S��Z����A�]fD��h��������o�����d|ǔT1���H�7p���b^����_���$��SS�$;��,���v��ɤ��G/s�=;��t���,�<zVP>=�J��Z~������1{�yܻ�4�VyGւ�|"�J��lqo�� ���.��Ü'�Տ�ֹ����]�h�i�������4{�Dp8�Z�<]b���.{y��1j�����F(��T4O�d�3u���s���%w/��L��ֳ����[u�\x�����m��*���C�pYp4��gB��](�B�?�t��C�y5%6���0��чt���a����db�QgT<F-�쮍58ii[�&����o��H?;ĪE$����TX�73����l��ɴ�W�V쁪�����O�|����:�6j#�V����4�Q��9�{�j%S��Vl܉=�(��j_|�x�VO�P�G�feK�_MGy�q\��3o�.���"����Q[��j+q�W���ZU�S�	�^��M�"ի��{�T�c�3��������	sKn��%�BP����+{.�	��4�ύD�L�<���CΕ`x��^����Jr�};��reIƄwO@��{6�v�R�G���-��>���*6#��u�c�=��c {�̈Ǎ=���}u��Խ�z�����tͭy���t�׌�ߒ{�T����,��kW�����T���C�aIIg�Z��s�$[X�b��tv*+�qB"M<ͯ����V,�OTfK~ݻޟ��z��N�ŊE�CJpe��(�̱�/HL�O������O'�[/.��҆���+h���nqOav�#a��rۍo�zgg�MMz<Ή������e�(w���4���UT$�Z9�nʾ�C�Gk��:*vRC�/��n�?aR=���>s�����1pS������ݕ��<�g������;	�rm��%,���K*	���J��mX*�w�Rǂ^�q�����R޸�{�<EH�H�����7�[s;Kh�tW�?q�O��C��'G�W���Sy�t�k�z>lq�A����Yk����,�]�)�\�1��D���z4�%N�$���m�m�$�A���x<8��m�Ɍ�ʔ	14�i�3���?��pp+w��碌@��X��t��\�{$��Q���wf���obΥJ�=Z�z�)�!�d���ѶB3C9��g�#ḡog��cd_S>��'��w���n��dvv� C�m��%=@���R5X%�ٕ����=9�E�ШV(��=�� ����+g�Sc�b��+��.���-a�x{y��.��ɟ�:��Qm�'r�#5=+�V��l�H�(���@�ѮԨ%��m�b���ߥf��W	䳦W64
eu,��Us�7/rsSc�WGƍ�����,8_4.�p��G�%҆��~��9��6>��,R %`���]N�V�F��HA`��Q�8��~s���ߝk۵�Ru��A��k���q1N����5ImX$hv\��uD��ԑV�_�2a�ۺ�I�Iw�32���L���x3��H6��������2ȣ[c���~ye���`Hp7󺣜q- =Ȓ9>s�zH�t6~&E˹.�%��Ҩ/c�U�E5V^D�a��u���N�K�7�Y������3�w9þ��ߔ�u���C���2w�c���]�fK�J��Dk�oV���n�i��v����g�I�춳��H[����<����2h��>����*_��r!��˜=�}��k���?�Lx>?r1w�A=�*f�]�i��+���?��Z�j-=�[��6[K�s�ۿ�'*$�{��J4���T�Hx�i��写��v;xs�G��3P�9l����+��C!���^G+�y��Q��!�2yZj0�M{��$�==Á� ��߁�T�&���|��kC����'��S����Tڸ��"^zjB��@��i�u u�$En5U���� "Pu2-o=��������g�j��M��*[�6���l`�Qj� �Cc��^��/�昑(�v��S�d2Q�U�wa���ϿjP�i�`��HÇ֍j��Q�G��fY�zZ�R�(-3��8�xX���tQ��B��k�{�U%�iq�7z��Bh��g
���o������k= �u�Qc��S��4�� �c�0AN�5W�� Yz5�g�T5h$���h4bq�d���1Z��%z��i.c�:�uC&���Dzz$�E�`�߾g���4�?�l��w�]�o�@���/fkeU�{�yL��['G�5`ԅBCӞ3�8a��,W��9�$0�W^	|3���E�7���8ػmX�����[��ڰ��'��e@@ ������3�,gf�dV[k�HQq���y��� �[g�A�l�XU����6�:��_�Pb�3��k�g��[���D��p��o�NlPU<ن��](;g̾a�g`<Ei,q��?c�� Y�م�V�@^e
Xy��Z* WZT�4�[�!~����O S({�po2�}��bD0��J��CO��Ae�laV�"�so�JBl��U"�%��b�-+�6%�/��j�\d�ӳ���t��3�����_����D��� �Yx�0˝��]	�R���m��R���᠒-��������w���V��yk��-o���Ox���ڊ��a��QU�E�'��oC(��v����RjB�v�?���#��x'�Wa�\mљ���e ,W1X�Y.彏�Y��I�f��XE��͞�tW��RgU]
*���|o����w��N��j�g�-�H�:���'���=�_W�MX�i��sת�ً1VQ\c).��K���[��rwm��_\�k�[D����$~}�������H}�3+�K't>�O��a=l������.=UyA�	Ya��tSt�R��Y�;W���[4�&ZՠǛ��)�	���cr�@ݻ?ݑ���ͯiX����$���=Y
���^�q�]c�����>7v�����y�Q�J7�E������?S�-�^���B���]�M,m+��F�+A��[�].N����ȯwIow|(�Di��@Ttt��ґ����:�+��=P�L$�H'�!����莧h��A^�۩�yս���/횑S�w�Q�R��bc Nʘ�3���P�j�rϒ"��X��R���?�s�h
Ι�Ӯ���[}�;)����5@���6�m��2�$����r�������z��Ǳ@���.E�Ai�IEB	)I�R�F:d��iF:��r�{�{��������7�f-����>{��y�9 �-�Ij�_����a� Z�f�4͉����[#�7��P;���;��:s,R���X���l V������~O��߷�����x.�l�&��9�����=;���JBݟ�7�V]�MD�Ql�ت�Ab`�̭-�7M�R��E�e�?.��v������`��\%��$iq�&h�|0��a��u�g�ڨ��9��T4���aK��`�����cqNx{U��[�ۚ>����?���&[1zQ�����h��A��I�V����D<b��_ ���e�� �1:�_���Z/&�)�u��2�!��������{��b���,&99��'��쭿{V:Ŭd���G��z�g�P�8������b��	�8Ku����q�Q�fc�ȉVq`�7�Ȫ^�>�4a�IV��l9��ut�B��Q��v(_��q���ܼAn^`'N�S��4��4��-����ku9�Ȳ�����S�p&1��*V�����J�V�Pkh�㟡��n��hۼ*e
��#_��UW��a*����3�0�еd��"�c�q�?"��Ā�6��x�:�3���'�q��A����X�ٕ��y�Zt[�hQX`7�[��nC\S�2��ە���N?��+Z!ۊ;$$@(�w�}�`R�X�Qj�;��=(�=:v��(�Q#FGk�a(�sjx��֢������HL65�I�-j5��N���̠�%J,����ϛ6r���ѡ�%^H�6�Mq�޼���1��6���H{Nɖ@U`��"���NL&|��2{�Y����G=�c�!^�S�F�<��(*�[re🡶���,��Q�����p}u�ͳ��N
�w�~|�ڋn�j���,�j�Np�*�S��o�KY��fS���u�T6�#w��wvܷ�I��ȑ�i(��Z�<�0�'��7l^M����]]�'�z2�O9h���\��0�k#d�R������fqUR�,j����ΆoT>���I�D�ƒAm4f��$�V9)��f�j�=��A�vo�Ǘ���O���5�Z��<�\¤�&z���/F��V��h��9��	�Ye��Q7,h�VreG��  2Z⇇�
q�_�
n����#��gf���'�P���hB@㝂�Ҟ��ő�X��Mݡ*�7v{�l����dY����WQ/����ɓ	V�����"�r����w]�O���;�J���v�L].������կ�2c���X
L�ťƄ���5���u謪��@��|0��B����?�T���7��
8��#����^`}�شN�8�a��'�����B���'#E�/vuJ~���+޼���hމ�IIv������e	U๕����a�ǍU�A�#L�&j���,:�<]#Z�HB��>_���y"/����m?M�I݉s�W�d�&Z�	EA�1��^�w�[d�w/m:�o'��Jl�G��o ��T�0ub2U�ٌ�6���B�P���Pm��T��H>�����i�`�SB7�"f1��M��,b�U�+�_�\G*Z'K:Sse=�0�S��l��˸V��5:���r���C%�+������hV�iND݆Dw�K��t�C=TU�E�(�!}�8�k��@[M�=��"��"���Z��T�dr���_9̿�C)ƫ	�5�9�����x�����ɻ�gs�%��!`�IN��9 <0x�~����s�oŏuD�Bύ��:����������.%��G��K���E���=]�0�b��FU\M����dj�7�qo�I�46l��z{vVr�m�jBC��؞Í�;��h�y��̔Dv�4��L��x�wc�V����d�0dX��z� �&��s	0��{~w� +]���Ҷ��������Sd���Yԯ�����E�>o­	-���K c�}� xd �V��'L������ŷj5X�������q�yk�TV���7����=K��X�L����p�U�D��P��g�~>��8��M�q���q��?GM�$5'�?��7�?'Qd�s���Γ<!��9����9��q�������~��E�9*"�y4��y^�9��X�o�>F.֭�nӛW�p#~m=�Ճ�5ޭ�m$��ͦ|�fX*�����P
b���Q�E>��)׈7VJ|�O֟5r �R�DY-���ah�6$�V��\�9�^��0X��,!/�� [� �I�nl�t���b	@f�����*m�s
JPP�xOO�xl��@fQ�G �̻Uo9�GrN5"_��P]!�G�,�;xhKU�z0kE���*/�-��]� �Sw�^��������q�����S?���+:	�[Q[���%mL����'ۛ��W7���lp����b�_!��i��H�U_�/�1\pX91�� ��̻�����o�'�ȴ�%[Ͳ�jy\<w*9��i��릦��P��?x����()�����A�A8[��}ۨ�P�=���xf'����.���>f� �0�,�Q&�����3��`�'02z.'�b["	�q7g��&o}�sV�Z�J�JW�Qb�*:��A/�����[K���:��n���vf�sദ��q���m�&yfQ�'��/{"��_ϻQ��#�d�'�.�ʘ;��)I�|�q�8���jG��A�2C�6�xz�Ǭn�/6���Tq��l��~Y,
���`p���s<|Y��4��/��p��Q\_�9�ԠJ��~�:Ҙ"�ԗZW�����\��Rn�M?�j\f�N��@��5�i�w���hw�C\���!���rM����,9��b�>c�S���O	h���m�7tWY�΅��T���0pH��	��b�s�mA���շ�|$K���A}����R.��uK�ʀc0�J����*��
i��t4Eq�� `�4�*����kc�X��T9MM���2��w|�����6���ۨ�4��l�(E|��|�Q�p��w��ab��ˆ[o��*9iͶEg�[u��>3!�'a���T���D}� �����āo�5ޫe��:f3�\H	��?QD�ɸ���Ccկ{��<M������� ��T�n0nBh�"��~	�~gc��Т����}]��NS�C9q�����[����Bڂ�������ӛ����	dS�Nv�c�ĉ�3ZƑ����<�tt�B���f�X��=������������Nb�Y�Flt�J=0�+w��#@�h}ON���I��i�A�.N����x�|�*sT�`�i]M]*�@ᚻaú:�Ƌ赡���ޢ��b���e`��> U1yN1�	QL��}��?���<8@��J.7 ُ�r�hH�P�����H�\�͈́Q��o�xbF/ب�����>��g�=��o�mfM#Y\�n��>� �!�ie��K7�5F�߄�cJ1�K1+����9����xZ���.I$uJO-]�b�ȮȠ��ǘc�!v�3uV��4nJ������'�[Op=Z�Ԋ���(��waD��{����/�W��MN^��jQ]����}5_`���Qf��\�1�}�̼Zc�ևM��s�M5��|��ߢ�B��4�1�{L�4eE:�TT�(r�h^�KQ�0���0���F�m����l�����|z.�m�Kʞl�_��]�_��r�T�.{��H�kq��u���07�b6%�(@(��C��%��kO�R#J�}�;�67��a|���1;���)�#��&�l��6�߽�\1+�$&'{�Q�T?/c��`.�� ��"aM�2�,E��ĸ@4/��(���0��UYcn)/�f�������,�'�&��~~�{ɫ�ǹ����Z���FO�*�����􌾭��[�zs�N[�4u/<��wG$�ߗ81�9`���gh�j�Z"��i*��� �M�ʁg"��\MF�9!�N�HG	 �d�m����Q穡�'�]b������4� ��|����髟���Ft��$��
>��S'��[+�JI$�a�v�����U2���k�����nn~�KU+���I� H���h(y_`vO�� P�ؕ��V�.؄R�5<(1B��@������0��t� f�?�?�݊�r��@?����ZIh\
�$T�h�ߛ��)Q UX���)�E������T�1(���͍#U]�)t������`@$�z32��1k8�c��Gzq�Kߣ�0��b��#���ƹZ�>o9w]ii�F��8$ܞ���<�)q����5)']�y�u=A\7~�t�6[#�,�Q��v���u('A�s+)~�&j�Z@����=̇ޅ�'vtts6�шNC��Z�b�9��zu�G6��|W�f�z�hN��^ڐ�O��e�F�s97�gH%��:�?���Ǌ�i�V�TW�`��"Z�:��c�r�A�v4��,߁~�i�<�-g����lo�x���0��-:ij,��3n���#�/�G1���DPK�� K+������p0���>��a���f���^���/K��yR�
�z�2PLJ7k���2�\�MY�ԧ�1�G50��U�{����4Z���V�M/�;��&V��J��M��gݤ�S�l�t�s�xeL�C�Y>m礴;:�����fͥ3����� d��9}��w�7��坼�b]ыm����y����.V��V�&oϗru&���]��"r�w��=�gR������;���}ȃϬ�~w}��7 [$niOK-�Sբ��4ɻ1zG��]�b��7x�Ž�y��L�����G�����01S4kg���Y��/��q�N���?� 8dx+��^��-�{<���n�����oeaF�6��ۍ�7�����-Ƈ��}|?��\����n�ږ�h�YJ��x��B|$�~�ҵ�uMT��8Bީ�<���57�^yQX!jI5��pIx�j77����_�0�&��FM�XS팧,uC�:;��Lm#=��ބ"fS����s *�@aˠ���w����u_'h1�=q	sDA���� m�k}�_�pÝE�t�#��j601�F&�(I�~. ��g�9���e���z9�8�ٷ@�h'��S�	W�2�ă/e���D�%i^�����o��%K1�����?�b�� ���� Zuy�~�Ƽ>zv�=�'؎��;O������K�u�������]�p̐��z,�ѓ>�	7`Wn��b�ЧML��*���\��'���A/-N��}�	mx��V�6�)�K��ŃEr�&��l&�K���J������~��3fE󘕔x�^zT�E�-�AO�ߓ~FC?^�\R�H�����|UOr���~T�3�h��6�+�jxѽ�U�����@��8�B��6�,��3�Ɵ��v��H��xn'�JB�O�'�Ę��9%�p�����m�����#j����a��I��Q�@�
�t�[�Q��J�B�V`�Tc:i�H�k����Ȋ�Ut�]�6w��fP�6(L%x��"[��.�nxOꙡ��x�L)#z_��J@z�"��o3����y�N|=4����6#�-Y1h���-Ɖ�����S����y�$U��N8Յwd�w�����Wt!��d��7X������85���TrȦ�SC�OFurw�\/���º��j��䐊e@I]w^b�L`�J5:,b{KE�w�5��Ou���=�Ŀ�hױ[��q~)N[H���$��&mD{����'L�ml��>#�-ٝ��T�-s��&�imhV��/q���y6U���P&If�-W��y����1+�c�"��v��͇'o[<�Q�D��j X�n.�ޫ���;j���R�y\�������bo͡i<�㙙�5D�IfUý������_{��g&�8�OܺǱ����8�֣0*�m�1 �<��M6Hn{��mm�h�S�ng���3�M�臚%�MSP�y,��JV���a�kEl�E��R�s�NZ�	,��U�Tr���:e'lЉ��9Q��%
6�r����AuT_>Z��y�SmX+�k�H�#�ٗ'�t�PB��kr���9����MGG����w�f�~�����������g�'��8��x؍'l2�S�ѭ�1N�9q��輮��6���<����N��R�鈴�貨�[$��1<q���If_2�d ��z��l�I_���r�
bw��;|8�^�����m^{�
�MI|譮���tmM==+��� ���J�n]��F�Zy�ƥy@:1Mr����v)���<�ml�D��љM��^��5����B�[}�\#��,��������S�^5L6=�)�
'�ɜ'm*&\1|��ik4&�ְ;s
Us�{�������sM.TN4�?p3���>ps��vm�F�����ܓ���ֻ�X����h�(z���r�q��r?�-h:���u����e�r�h�'{�x��W�b�5bD?x�yvݕ���7����6���r��r�C�w�
} �<
�}��M�3���r{�����~�i���T��D��5�5Y��(�·ר���Ȉ���H��8�V��Ό����"T��Dc�1���2�M\B~�:��Wkir2@���zz� �^Ao���m��D�;�qX2�� ���1U[cw#��;χ��:8C�9Fl[�7t��	�N@��Z� �ߒ��y<c-�l��%��5cR�#�L���'�`��9-���8�	��

A�D�X?�9���o��z"�H��v�Y��;�r1T)����x�s������ϻ¯�c�����3�qF'����֦ㄪ	x����Hp����n�]KTo{�`��h�|Tdj�}"��|6@9;H|����r2���9�F�����5������w�����1�~� 8���~�!�Δ��h��9۽�+rz�������~���Kѽ�G���s,�e�Q@,gݝc˵̯�u0yQ �j)ʺ�mZ��3����Mg�o9����+1����O��C�����H��i쬌�,����Ha�.6i���M����W���Q
��) /']1uC�^�v:�狜����R�6L�/}5��V�걠K̩�`Ô�	�C�|�����fy�6!?��zjV���oe&���އQߋ�G�g�1�@Ϩ��[S�Lʡ�ۑf��p��V��@�b�)�RQ�fY/gn�I�[�^�c]�o��Ɉ@9�"߳^���SQT`�@��͏'-Z\�����Na�&�iV�d�t:�<�X�O���:����z�܎�c�7#e��(��D�Z�7]�^E!�(U%�k�]�����^�2k���L��݂J�~���d�N�&e4߼��e���	d��&z*�,�.;��;���K	�v��T��H� A�_���Y��m~�S����%ߢ\�w1=׫���9[P�0����_F�;�;�¯���V�fsY8hޕK_W�N��iy8����iEl���m#�	cgg`A����"���(߲��[>��~P���$����5Z��x�rDn�:�$�O#pz\�͞�=^�'v"P �,��W�?��Ǵ�o����Ы�xٕd�w���vn�?K��nc,K~�U��9˸���Ǵy��(�
2�W���:a���ɉD���^��k�?�r��Z��A����>�fi�������f�װ%���@.3���հ�[�)����:�>7LX��!�Wy�h����Ф�����WG�܋�� �g��l���|ܿل�I��|��������%���|�e�9��җ[N&�܂�	馻C�<@S�(^�y5�+2Pe/3ԟ�3�"��B��Sˤ&KȞX�cz\_����N>���p�Q��ɞ\sӮd6��6���-�/S
�4�2A~�v�_����*L��{�pT)%r���c �Է_�x(d�����a�لQ����Ozuub�9w���L����,iz=U	��Ͷ��x�B��08
���Ezs�s�����q=|�/�T�� O@��`t�"�y1����x��iqJ��Go�pz#�|��y8F~�JE�X�j��|�S��x{	���M����R�Q�<�f��9p���NS��J:FڻKKo����궏�D<g�{�ތZh�i�����ܐMZ�[�b�bmI����6��q����!7��k��n�߹��Pr����3-NvswX<�V�������V_�~�g�U�r����-��/W��S�`�M%y��}YnL���-��J��Ř93g�����"��89��B�I|�]\���Ʃ:�C|��D=VǍ�T���D�������7�2�j�$���ظ�$�:m��?z��#�.���~�B�gyު�Hh���=`{>��;�w�}��p..�����������i�������G�Q'٢�t�W�Х��>����Ŝ��ϋM�����'cD�'�SI�W&�]��p�f/��������iEw�a�?|��!�i4̞xkg%�2[p�aC�9f!�i��m��`*}��BQȂ�ݸ����
��~�B�e�YCD%�o����={V��E�2C�QuW�y��s�$������ٛX���G��^K=sȟw��⬝�Vf�Qo}Tc�x���ˏޕ��[�ߥ��%�?��~F&�>O��9I��U�HYVo1�Y�z�_|:���'T饕U߱���ϱ�&��|�v!�(/�G鏦IG��ŉ���u��m���zu\�~�{Ѡ��Q���ǯڍ}HBY	�����Q,�N�#6�G��L����C�<�����k�Rͣ� �ȭ��	9��1�r�i�G� ���-63�5�BBiB��ת�5G��^�"	�c�ܸ�~��C�k��.�^��U4�c�A���f���� v�d�(cw�ۢ��v�V��᠑���4O I����r4���2%&��%|*�?�MqΊ|���y8�G�]_`��K�K꿎��w�@�vN���]�Y��R�����hoa���YV?�T=�K�>/$�/Ù��ɔ��v@	�j�Ps�㙙�W_w~��B5!`o�U�����ʆ[�W��l��'>�3�K�D>N������sD��oUi�L,�����a���Kۿf�p�P(�dW�|S���AV4��ŀ�pV���Z��fO����H��E���J�v?m��^0�M6"�"T��*��6��%�$ �H�?�$���h[��,c�(�i8O%)^���͸�gXE��8�v@UGy-�~�V�y���&7�4�-U�����r$c�=�����?n�\)ɗ�<y�G5�ZI��c��[��0g���n�����r�z�H����(I�5��+F6�����fL�{�6��ȥ3;�&���S|9u�n2�Yy[]�y)I��1�F�O�7�o��O�t�&q���_���T��� �m�5֭�t�f��u��ȳ�?J��b��%9����CՋ�#���F��d�O 7z��~��3l&H�%��L,��̈�{^ȿ��s}KZ����һ㏃�c�e�-��&!}�W�'	�[�}I�u�>ú2i�=S��Y��:,my�=-�V�c�d�&��%�BT^����.���<1~@>�0��7�V�S�[`���vQ���.x0��g"B����#�)��
������T?-�*�?w�ut��L�Q�6ʕ'OԾ��|myjg;�vv^!U�h���nr��x��_���է�V�
�����N�o�d�G�e���O���9IdW�+}�rsT���M��q�
�yY^�Y��n�ˏ�ik�_|�-������JZ�z��×x�{���R�E���\%؉7���0�҄%c
�&�Mby��3];��O���XX��_�k�3��C�_�o��Ng��K�/q��d���yDr�r�P�w�MR�{�+���w�y/ݹ}r�O��js}��[�����eޠ+�vB(���Gx&|V^8�dX�T�P'�E�����M�0�Z�
�U¼uN���� �&w���M�$-�{K�z�[��iiߘ��Sr.����{�p�]؅�[ͽ��%1ߊ�ӱ!|��r:3�T������d{c�1�-yY���6��EQ�L�S�(O��h�]e��P	T��׶��ӛ��*�ʾ.+��#�t���`U�����F��[̯�Y`��5$�����~�E�{�ho~ >9�Rs�P� ��X
k�m�����DSv!��~I&�
	?���eܥ��Q���;���ƥk���VĪ;L���!q�������E�gV"Y�>�>\؝�+A7�m��c�(r���N���
7��!���%\.�<(�R����r �A,�*��C<�ϣf2䈙�,gf���r�[�IJ:HnT)Ʌ{��E�D �Ő��27>"X�j�6yYN�y!�@W��Ȗ����#ܕ$�(}�6O��e^�rԞ�z��^�D�c4�:L�t��� \�l]5n5�>E�o�iB�p7^��&��&�u�êby��ѓt�� �ͣW��# �����ȷmM�+jI�Q�(C�>+�lgf���u�f��(*KsR�_^yA}j��;��}}k��u����$jB'r̔�g��|[A�J�9�6�?�؍��*b�.���1���$��$<����2�i�ՒS�d���rN\�Nugi��'[���wށk�S��tzu{ �m���/�k��>�d�\��^��!=�൵�`��'���d��Z]Y�_�Ժ�[o��}5�S��#�)����H��`��8`c*4b��|����1�}{��].��Z���#��퐪��)1��z�?Vױf�K�|D`�K9�V:6��Df��o���}�b��6��5S�ȅ�~�s�Wb�$���q�¨�BSS�����W\����X�;��[��wX�Ωuo���8�a�¬G�;�A����d�v]2��9Ju�)�~�A?�b��S�6+�RqH�5���
��Q�>�
|6Z�Å��
�z���	òq�>"�w��0�p����:O�Q�R�/�ll�nG1\q�c{6�U�&��1���V�%{�q�L��y�5*��&�G��y�,��Z�M���C¾,C����~#�`m�[�C��߃c�[�V��i|k�m���y:�j��v7�i����gI^Je�(	n&,)X6����<�o��Fy�;�$�NNO��΍r>rt5ͩ%�V�T�|��=�4��d���C�{�O�����0�]��O���Aa���8�_���H�Kl������ֆC�_��R"�R\��p@���3=���N���I$S�s'�.����2�/ ����L_�>�1
(6�w�;TH؝�=6}��<'�Ē��rT mj˾F�:��[a�)k�3j_XVM2{ؔ���-{^Ha�LL{�fΖ�Ő ��U##���ѝcr�O�p)��g#�<�=�"d�������{�?�ǹ$^ύ�l��~E�G�����mm�����?#킛�AFePH8r�f�f�-wG��[xM1�̅�x����<!�d�;��%����v�H��麪�	.����C�bD�L�ԧ֋k��b���5g�2;{w�A�
ۚ9yy�&&&'�kk��i���}��P'߼�w馟�O�z}Np}��i {�����AZS����|�SW%�h��x�˗��<����{6:���nsb�5�JvT��Ųq+[a���$�L<��'
�V��W_	mI�oZ���d�\���^�9p�����#��?�I����u�2T�Q}*�!aU���y��������G���/�w�F���a�U���[��_<��6���u�m^>������ޜ�|)�>��Ҥ��Ȍ���_�g1<]K�)�A�����}�Bdy2�GYYY�a�Q
x���������ce��gB���K�����=b	�).��5�z���(�2V3-���s��\���P����ڿuv�k�h��M����q�-)���8��!��a�O� ���ͪ58 m�� ɶ�u=p�4��vnu���~�G|�"�<�?�T@�'!��݈��5SE�S�2�&��K�����Oe��H��/Ï���캹�z�/Z"�4�_����L2NEE�������G~��{o����k�-4ב�a�-,���j�T/�0X�D+�W��O6�=x��[Yt-�
JH�2/5!��٘i��sޖ�aV�`b��O�����K!��d hn��ş�
��%�%�V8D���;��F|N���p����Uc��_�Fy��9	v]5@������m�w���#�N�u�*I?�SܷY�$+H��Þ7(>te:d@�;��x��A��M⼐�T�'�j�r�0�E�.#i�΂���O��)��F��xٞ#�~�N�H�_m�${R%h����^��=���g j�a�a�4�؅��bHc��{�ۧ�f��ك&��� �χFF�ǌi�nc��"��Ӂo&+_�����Ud�G�Pg�c�dg^X��9d0�Z�=Kkg�;�߻|A��Ҩp����'G��@���w��RU�lWU �Aȳ�S���`�;,�X��[7�m4��'���w7=�/
�7iP��5�R1��-O�V����w"Ք��S�nM�?S�K=�?�!-T�*�#�\�S=�wf���^F�9]���|T���k!|Oy�f�����[�暽p�N���[:�\��%3��i�8��$�-)^Jp1)�N��C�����y�=�b� ��6HY(C�z辶�5��}Ն���p��7��0V뎹GN���xn�D��3�^H�٦�m���f��z���.Ei6�}���'"�
AYO��W�p��Ԫ+���������v��K7Kn��*���_�£ׯ�'�L�5��gv���Y�$����P��P���Y}���w�z>�7	�Zm�Ql�n��D������@��m��yQ1$)r�	��iS�m���9� do�f�5��/V����chȊ��w�Ą8��}.����@�������6����-�4�)�eh8�� ����}�'.q|��]em�Y�T��k�5�'-�ؕ=Hf�ȕ�3j�R��_�/g�딾�J6��#I�}�@��d����p�y�K�wq}������j�g1��k����A$b��$��0D��ȈVye�|O�e, ��6ާT(�7�L���������2$2�����W�? �8*n�
}�u�@�%���'��b�����H�j��G<�
�J�������o�D���r��1�z	��x��,�(+ߐ��;�`{����t���a�s����g1�c�+7��;w��WH����ݮ�A���A��𮡜�h�[0��		x>�5�f��v�K�D���~�g���d kw�o�
�Y��wܬ���m�}Z�)���+-�X۴i�>��G�z�/'5$��E�v{>m�[r��j8�*6ۓ�M>z),pteZSgw�z��˵�%O�{� p�R���į4ֶn��d�'�v��������I��dݛBYP���-9t+�K��~X>dV �6� �1������Eڐ��Q�/�/��hia���EuFs�6�ttt\/(��@�5�/~�E�sA�d%�B�^j`pp���6�P�����Az�래a�> l�V��	�um���/�k�>u/_�UK��YL�	���H�m�5^�Q��7��q����K�S�$�ϝ-H��M������N�ǙE�k�7"�u����ȕ뎓����J�
\�9�x�E0s�5���UQV�m���ꕳ�Gm�#(
�-I��A��o��eݬT��a<z��1����%o���p��sh�w ���6t�{FF��G����$��i����w�ES[�5�{�b�:��;E
��V�����-�J��G���y�`�I^,i*� �� 2���3T\��Dy����OX>���eH���A����[J�`="`:s��)��q+��r��,���Q�W���i|P8�0՝;�#l����-.�N�u\���'��ld	4����եߋ�s+h��x�ro"b�}�e���@������Z�Nc"oJ���A�7��_�����0���[���1���_L!/��Y�MGH�	��䛳� ��Q"��vdo�{�h����$u�Q�@.|_x%��W�q�{w�qN�I~�hM�1����O���d2�r����C����A��M���Jb[41~:F�T���R�i$�Td�����=(�`)��{�
��G����\�]T�:@�����r��^����aPY�LͲ�c�އ�����<�}<<t*xQC����#�!���r<:\Rc��;W,*����X?X�x���<�Pc%.�r�]�F�;^�.�Ǒx��b=}77]�U�y���
n������'�Ӱ�wx�R'؟؋�h���vc�f��Q<����	!fn4`c5̑�$��ʳ��id�$Wɖz��^m]�p(w�GX�\\@�1��b��k�7��MuB�hZ��_qcأ����e��>Qm�DiL�������f��L���=UL �N|�4RgV�������`�8���Ʈ�K+��/y_��7޷{�A՚�����e�:'Eg�ϑ)��"��S��>�tYt`x�"0j�!?-�����V����@�HǄ��x�s�S�ٽH�����4�#2��m��:��j$�J��L��L�oݽ�����"�v��� O+�Դ��My�ɦ���|\�v���q��b�x"��FtW���nA<�7�4��^��]�N�ߨ�(�Ҵ�I��������wn�̧6i�i�pu�.��M�V��I`P�08��H��>�(2+|>��=���;��7��n���N��8[��,�:��ੲ�M����2�6W�g�X�j� ܬ�C���Z�b�s�ъ!��g{ko�����";$r�?�f ~��\�6�u*�JSSS�ƞqbr�İŧ �j�<=BT��U�thb��N���ņN�#�����GL
?ˋ����t�W=/�:n���Ȫ B(7����7���a_�W��&�06�c�p,Ҫ�Za���v��oF}���
�Lqw���)�:2�QZ��9:6�_[[{�`L�~1�,�K?�tw��&AymdB�cfd��R�S���pݦgN�?�x7��P�~�Ɓ+d?�ɥf�|ڂU�}1����SY����5���턦�������W��f�F�jFx����!����tL�G��W�*�PavB�Ѿ�{�U�g��d�(���Svf��n*����뽫ч���F�-O�ǆ! KtKt�n��/M�/�~կ\��#�<����y9��n�f�~��M_�P�η��~oL\ϸ�߫?ݪ�f��v������%��	�d#��I�ɛ��1!MV6�>�Iyԙ�8n蔼�VdV��
$^5��G��������n:!jp������+�r���'��I|����RK�O)�2��>[�4ҼE/���)W�/���}���2�L��
¢
x����]O��8�Pm��Ɏ�\�J��P�8R��S��bp��Kx�^�=^S���6���?j2[�D��Y�eˑ����Q%��_�����g�'��y@)1������6
��xT�x��ݱ~�D/�	��KjW�Rzܻ$��J���j���(�yg$c�n;��Bf��'��1���s�ͦe-��T���8׽�S��������H�gc���5��I_S	a�K<���e(���T�"�{�=?8?�k��G�Ee��,�rI
f�lm��Q�d�;��~���+F���ƪ�Z5|]�N+.��2\A��e|K;�K� w�r.���C��<�a?~SHI�W�Sp}$�J/����p.u�,C�fW*Z;i�(�{���p��ȳ�-K�&��� .��)[>==�FH�u�h%"c��$����y����-yړ�-�@[�k���=�oiy��sf������y�-�z�=:~��:㱧\,JN��;�/�WQQ�sz��CЦ���`��3����{����#Ň>L�{�f<y���_q�����3�x)O��[<I@�D}�z_�4��w����;���[H}�U�.�ۼP�}5e��wjX��&�1#+,DG���ڄK�d��2�ζx�1L��%]����������q����z~�a�R�1;���}��ϩh�Df?}n�����Q':�v��R��)"��p.�q1i�	ͩ��b�J���&N���D	�M![�����~���L�t���a\pZ�h������{���D���!x"�+Ap�(�pY�<�e���<y�dd����9�	�l7���=4U�e@h����#��w��DSs���df^qژE;��YY}��r���u_IL���a�g}q�E���#R%������}8�F�g��|�W����4�ЁbU^̜azf��X��苷Dw���OE�ʏPG�����#�'�v���O�����e�v�2w�����G�ҫ�t����Y�Tf�:MY(uq�<jr�tG��$΂�}��he���f�\��v.�+eK��Ǎ��Tu�G�Q�Oyq�fIC�(�L��x�o,���)��x RA�ٷ���RU��$�^�Hr� pD,���}�%�[�(0w�+p��,f��3^pӪm��E��^M����J]���ݏ�w�Z�ͫo���)C�ٵ
0u�����]�4���~>��A><<<Vb��p�Ly˄��|�t8 ��ՑlG�Rin0������)%�uB-(���ב���#���t��Ru�|���+L�1;��h�ӪaCRg����뫴^����wno2�P�V���MI��k���8�q�"�N��u��sb��bp�}4������yv�}L�$�[��'��O5o.��z��R���65RhYӒѮ|���~2"�o�\h�_>P�_���i[���2�p�\��@��b "�MJ�� ��jU��s��P	�(Y�ʏ�M�)��)���]{1����ڹ��J.M;�7o�c_�X�`_'����Pޛ�&�u񥮎*==ݟ��R�hz}�m@Q0EUWW����/P3�s�p\^��Y[�Y��A��Q
2&H��� (T-�)+9ާ�TB�����SQ��j��~33�G�������1�,����;l��ᛓ�ׇB�~�Ҩ�͗�+�WP��y/��v����Y#�5�.���Ol��Ll�ҡ;B�,2G��܆C�%�0��f���6������S�	/�;CY89Sm���>+�T���'q]R'r�R�$�o�}��[",�s��� }�����U��;���w^�E,p��HuHF�ܲ��+ϸ赁�F�ߢ����<pJ���m�83)��l�9C�]��Y�L�@[I`R�w�uk'��pe��z�E�ϭ��Qb�~+[z_9�癭�?������>���"!�"H��J���-!�ҍHwKH�t��đ.��Н����{���ُ�zԳb�9�kͽ��ח�!����V����&��}�v8T��Rr[/ϴ��f �������]>k�mAro�@Y��IO�f|�L��x�c����s��\��č����Ɲޙ������
��L�oW�{'���2an��ܝ^��XQ����@��ի�I�0=�$hu|qe��
GFN����>��Ņ;;;[�T�=>s�H���7w���P93yId�AB.��9&�_G(�3P�!!X�dX_�*��|s8T���W�N6$<��L��������4�@��N�=NW~�𹽿�Ә��X{#���'�����͟d%��~��	[���R)2/�P֎�Uib��ob
9z�Aٹ���\k���;9���8���׍Π�����n�`���&=���O!��v.�U^ẫm�!v�w�Ls�q��,l����FM�1�w ���@Q2yab5�oo�iݔMRI�r�}�3��'�f%�U�'&N���u- C���3���<�XJ�ڵr��;1����굧�Ѕ�>t}�������퇯#K��P��@�F��Kh�dߥ0���fs��Oɥ#�5*�f%�L�Ϙ&�|�����y��_�F�#��݀������e._H4�Qt���
~~�N�v���?��#��%�w���g�%$)u��3%.Җ���@�>�2�@��ǀdIBBB)e�{��~��e�-�-%-�ee�J�&�%5ޒQ�&R�>0�����ru��_\^�Dw8���h́��>��\�z��U�"�oL�ޘ(����s��&"m�F�v�/LZa/輏"L��ƆzB���11�
�O�ϥޢ�ƚ8y��H�|u�r8d�Z{F�������ؼg���'�S�[�J���m�ɷi:�<z����wJ�@̱���$�v�����u0g�wg�(���d�Eȋ�(CF|�<��Ȝ#pK�.�?�[������(뭟��Ò�b;��I��8�4��YC`� �F��� y�椻or<�LyĶ������X�H<A9�B,	�b��of��߽ٮ����{�E�d�[���վ�����s�׷{�>� E�Nm5ʞ�b����X�`��U=2��J��o�gd_~��}T�k�B�y	�H��R��Q/jy�Szv�G�_�P��"l��cض���/�{#@�e�E
� �{�>M��[��v�`<# 䖺����[l�@s����he}����P�f�7QCwߟr=8މ�{�p�S���;����+�Y�o���F8"������F}w��3��(�I����H��S���MR�-�,Y�P�h<}�ڮ3����8��}>�s��xG���Pkzz쌡Ȉ�����|�t���������n�CE_D|�ˠ��0�HE�u����$�>z2RJ4��bX���jd[����ǝ{�=wC'�����JlP���AZ}W�����E�i�ǔ�B��ժ��� 5�J�6i̓�b�,w�W��.k�><�U�pj���7�B<R�ጿ) DMMMw�����Hd@ɗ�`[�P�[|bo���g��F�?� ��`�������FZPwD�}��m�pm��WzǄ����DPP�߻w-�����1���>�
���Ύ�q�5x��֣��D����"ы�i������p'��s�a��#��,~�P���f������)�%H�5)���ޮ�ܨ˜\UE�H��>j�޺��>>M7���rX/j�d��e��7�x=.�V߆��J�7O�A"�޶����tqqQj'�4�� <�2)����Ν;l���,�&��x��tyKC��0������]�?\�8̌��r>F4�Ӭ-�H�Y>Ackkk���5x$�j`]�X�M{b0|""Q��`@)����00R�����ݿu�Z�/T�b�aaZ��W�y������Y�=W�[0�v�lSz�_�ZL�].F���1j��0H'��::���T�����d��������Z%/�?�\���e�৑�U��U���9���B�f9��}K��?Q���c>��z�����p����7��@�Q*۸��(��������B����A-=}}�@s�@�P]=��X��oy���9S:�1�ߢ�ˀ�l1���Xd����x " �/}: 聓����B|G''�хg�dd��Id>c��]�����j�L����k��.�iK܄Y�Ӡ�ِQ)��o�����m!w��wD��rpPj��f��P$�3R߽	xRz��H1k4�ߠ.�h>!�'��P�e���:�]��M��5�;�o������.�A)�^	C�6�����<ߔ��W�iyG��=�=S4�3เ�n�ˑ��G�0���XqG�VF��R6,��G�.��X��0;����Բ���i���f��7`�u�M˜������[��)�g��xcĴ��`�A�o{j++	&��7�}i7y���(�q��$N�!�RPP�n��D]D �ϽD���"51����C�bbbr����f;�ԯ���*V��.�	�����X��������r25��;hfL���v1����i,����Y9��8�O���0Hw��_�� ''װ��8�������f���"`����t*%wy�z�6֪�g
[H�66,�yn�0��a�^�i�FA��|tt4�i/b��>��|��w
��jA��,��>����)����1!ǃ؋�����|�*(���}�ؼ~�ĕ�K�ϳM��^�Ǒ��0qOL�O�w'���&����w?� D�T���%9��-�F��G >����߃��0_�b���� �gb�c��.�7H�1`500x-.�����+k�xu��U����{����ρ5���'����Q
?�咈�J�NG�ﱿ@�~Y��@WqYb*=a"~sũ�Yy��w�:� ���&�8@������c�7c9�T �ѽ�{(*'��<�Rw�g!'����uy�(���ej��^l�������5gG+��$����^B	��s��)����\-��e,�������Q��uH�����@�c:��`aQ�!�|<���>���e�s��)�T��Jnl���h���񝬬����yZ�9 !�YY�>p����������@��@�zUK�p_^^�ַ4eUiф�j���/>L�����7��c~�yI͢���?0%� _�8j��z������`���;H�\���DX=b�X	;>���<���; �f~�&ce8?�Z|�Xcy�e������>y�Qq0�o9b������l�d����V��QdH21�`Ee + �h@�� ��IZw_8:u��<_R�4a��M��Ұ��m2R����uQgA�z�&�ņc- n����W��Џ��U��{r�e��S�c�!��X=�k�Oo����|ҶQ��/��*u����ycu��(j.����B�����AxC���1y	Ւ���M>����_G���i&0<�����C#���Nŗ3�=^e�Tj���tݍ���b���$2������x��
�<��
2-�*���lox��z�(5'5D�V(��V��֗��EG�W1����m��Дs&H�Y6��)]��G)��g�?�J�'������6v�!h$�̼</06�u��	v�H�\݆���"CM�|�Y}�.C͟*�k�2M�Z(4��4/0PO�W���
ƎQ?6��<`PdT��A�4�>U/�����:,���v��1��7s�=���~(&��활*,,��#��M��_.%T��R���Cו�"wk���p�~�@s
�l�H��� �W��m3eu�.���)!�F�N�ޱʑO�=Z�4�[R>�X�_��5��tDZ9��,����ga;�� ӗ�}�9;'N�K4?����OǇ& ��1BĞ�t��xzz������r�h�.T,$:113��u�~+	~a]�+�6\W�τ��?���.��~@ $���ڍ�Sd��J�,Y&r�Rڰn���ŵ`#�'%����������(5	�J�^�F�Je&k��cn��ǈry!ɫWB��ˆ^�%qv/�{��A�&d���Q0�8��= t��Nw��(�mm��)X�;FE�YyjY�K�/�)K ,%�I�>(ۇ�Q��de=��U�S8Y�?�U�S�:^�?������W-p����z���>c��Qxz0�.w��^�4vU&����H��	�����{=`&��ʣ""�KKq�ѕc�y4j���	�(1�Hf��vO7�~��َ9��*UZ�=�}p��`ra���������]�i�_1F��i �-m�I�</YY?766�"#9e���7,Y��<���P��38��(&�����P���M��M���6�k��s��}@������%�eC��αo��Y1g�������:�
:��
�n�F�j,Q������ E���$Q2��azs_J^��B)o0w��b��}W"�����Ì��*Ԏ����W�z��	
��h�#-�9.�>��م���l�q
m*c�+y` �a�<����V$| �`}��MF.3��`(�7`�n�bs����.Ƕ���� ��Om)���z��Y�K�&���4�O.��txr��eP�t�1@�6f�')!��(� p!��B�Pʷ��)|?FLq�^�������bl�a�U�6ݟzQ���xӉNk�St�/A�	?ොq�g�?�5������k���G���5 h�a(�izF>�>g���>8��?0P8&!�  !!a�ؘsC���_�D�����Ȱ\�R`���	����-���U�V�(j
��|c1��9��m��{a<85g�ݷ���OL�+_���N�[7 ى~eN��C1���н�?`p����G���p��M�H=�¦U͛��E��~��C���� �e������5K�X>�U��C:�G� / 5b�ajJk�U��2EEE}��b�͢�=��ꠊ�J P@ ���qC��!��Q����b���n��p(s��bN��멙l�WD�(=rt��Y�^��V�]��s��w=�/��� 芑�?����IW�h�_��	&��}���{�S`����Ot�⺇.�tѻ,�w^V��EY��<�;F�L ����#���;�;��֏C�t�sz.��YY-�8{Р5��nw���k�Aƥ*5۝���sQ7`����7��K�o�Q\A�2�
�~���{��-1B���F|Y���S;��~�C�_?J�yt�Hq
j�S<5س�&��_����{���Ǌ�O����ȅ�JJ�g>�����Jr�
��V�Y�S �AG�y�ݽ	�w�N��'T��f��cu��$��Ey�+/,� ����OK����(Pݕ�+o��d9�DTD���uS>����I{�Iz"��H�&�TҒY(���d8�*�\�"yjNz��-"\�sk�9��E8:�O��E�`�s|���ԅ	V�NY����,�m��?cK�`�QX�ڒUu-�Iܿ(w
`���}3�g6�^��}��U�	��h�^L{1�xף%�7^�yV~\�iD~���6$|�fT�����J���}�[�y�5�� ��O�f�-�%a�wv%T�Bf�_U�I�j���Ė���a�����
A���~XU7k7����ZW���� @W�#�x� ^�S�`	�z�>))�(Hk����ӧ�� ����L�핿/TB!���0��H�L4d6��	��i �V5��<�Zq@�%G3����xϰ�r��9x\f6��ȕ��W�ߣ4n-aU�r��+�}��q3ff�o��n���j7�����4f;j
&՝������o�O��UU~���A�E��c��˿�/+9�i��'�#����ӗ. ȗF��O�+)��_�V(���=��-/O��E�y����UT�Ć#Z�?���~`#� ����(x5�F3?�xBvp��@� 8�x�xV�� �#*@0!���d
Y�P���*�<�SU��4�̗�D�hR�U��W���v������g,��;�K�#Z�d��s�Y���^:r�{O���^�/Ŭ��9U�HX=y-�}�q�Ipt��m��u��rJ�K�xq©B�ʐ�/�:�r[��f,;���TtYvJ���	D���f�ܮ#���΢���-s��F��no�b��b�y�ʺ8y�����g5�b����jdb޵Ї-ɕ,��=��ő�4�e���Ԝc����/\�NM�׎�~�Xw���?N�Ǌ��e����@j�t�Ç9��"�A-i��Ɔ�D�#C��:��ĖٞHz��u�����ݜ��b$��F^?#|Ѩ��Ja%����)��#���uU*�YŹ�<� ��@Ǖ]Y^�	jyG��iϤ#�[��=�kB�gaGs�z�2������������ǯC����pͳ"����˓ob���k�p�� ���')�_��������\8c�Zh��p�;i�@.� �����V��`�&�k��1�8hw��ƥg���n�ӆ�1�n�;�y�϶:���� ̭J�c��_C��@pyκ�_k�U�(bp�t|r��F��f�6///5p��9�׭���X�뵷��I�ۉ����W�Wh|�b9n6?���p̪;E�����}�/{��UޢK�L&��&r/�I��B�tw1�r�Z�u��>��T�ecc�@�_��˪�R��c67/p�
K�,+��U��(�⡅�|� <=�<�u�I����S�_�M���D�"W5]^�
k��Q0���i4������>�劙my��9+�r���	�:N{=,�'�4m�$�{Z2�Y<&}���X�������cƋ��ݳ�n����0?�|<y^ɨ� ���mbbB�E<�G�X�+�=>��6:x/mAMʐ��i?y)?Y2�I=r�I.e�B���lIN��Ą 0�ʥ��/�^@�߾���-�pn����t
��;E�_W9��@4��71�IK'/�ep�?h���cq.JS�9������.*Þ�#�d���V\���6d.���si��ۆa�R����c���jf����-��"��#PPQID�ie�A�S�lU��W�D}�����i<���kg�/ق��(��/�*�=s��ڮ�������B�"s���z�M��/:��ggS���m	Z��=]�|5����J�Er��2���>�u�S���ٍ¹H�����7+�\Ը-�B����j����˖rr���a�,.vK����� ��=?���, �z)+#qF��-6�2� ��8��-��>W^e]�=��h�b��w]�,�w�-}�8V�q������v+*
���>I�<��X+��������d_X��L��6�hf
G9�����ŉH2>W�E�w�\�sC���
وI-�� b�+ ���"x*+��9jftMT�Va���4>���tc�g�kW�V>��
��ֲF���C�(d<�a:jd` ńOl)fk[���)����D�=�/^(���vq�ǃ�x�+���}A^���ҥ�ei
;E��"�|K*�)��˻^�����R�zjQ�baa����,���o�܅i�����]\N��41�}�&0���Zɯ&n�t�^8��Ө������u�!H��cV��5["�ey�����о��?>�}e����w��T�/��'�C��-�rG���O�Zf�ΎVl �c�<:^$�w�X%7�l���y�k`�R���]O��1RZ5�J.�(QaRTTF{�H̳�����څ���^�ac���ngʑ�A�P%zib���qP���ά�Ĥ�~�%��R�N��?0���=�>ZLeF��@$IaR\\ �2f����	�Ň��AC�M�P�5�k��ui�iFԵ�����.����٧1JfI�Ne��3�*��J��s���~��ھ��VDY������O�H����Y9`����u%_���UTLg�{>#*��"�o\^L�t:1)�`$ @
���:9qI�� ��1����H�Pk�aSJ|U276�[)��_]5��헥������e(���ة����x���E+]@W����VT��0��E�3 Q7 ����1(n�o��QVj��/G�=@�&���}�/l�����6�Om�T[�țZ�W,� |
D/��7�J�k6��X�_� Hs�{�YF�%�o�����W�f��)8����r�^�� a�T��4ŕ�
¡�6�G���
W�Uۀ�D"�x�9+�,��)|�nUc���?,���4X�eU��䝜�
4�8�k����|����#xv����%0b_��І��y�j"����4
�L���RVV�xv���ӷ�$7�i{���
�N؈w�4Љ^�E_F�����e���m�Ћ6Z��7�F
rs�=1y��Փ��!�`A�����r��hFr_���nU퓘���{^�Vwl�0֔���426&�@��)y�3퇚2��vL>\��d��bBbs:,*Pƽ��������V���7�ǖ�B���E3������R=ǥ��_�ж~����!��m�Z�Ҳ2#--�_g������ �:3
�
�N�Ow5�Kњ�YY}��GfUK�\�G'�q������݌5Q�%?Yj�NC�@���*�񔍌����"�e�,��T��2�8D�K���w�ხv��㸼�f���=@d������:f��G���d�%X�22qwNA�v^A�$dwCì��u4I�K���[o��hH�ք���§`�\(���t�A�ոu�(B�)���XN���4���`b���Cȏ���G��H8mŠ���S�ת���N%Sh�ԯ���~�ӣ�޼��ap�I=�&sA�"���ĵ�CG�,��u�z2��)<�PV�]��IWU0�n�tS=�1���&m�.�E���U��������
��D3��t��HS
]��"�M���2=t�2�a�_���/����f�ꉳK�7[ld���;�ϖ��V_���5iv��Ә��x\��]NW4�c�$J�G4�^N��nl9�
@n�� �oĹ�5u�3�e:�U���=��k��w�B�2[���UnT��UpL�[���6��,�H署o檽��3N�ܠv��$���b�
��"т�9E�Gi�f�:��x��,$+�F�mk�Ҿ��WB=%�s����(x����[Ps������F�.3W���u������A͛i`�-S��4v���ȯ�V�ꡕh�"ٵ��F59�����]Xz�=W���VT�z�qxT�$�> ���^��7�v�\�bgU/��I�p?=�"��ʛ_r��n>8�$`�l����ez��O����?�&AH�7���0��vg��k(�j((G�U
H��+>bA �VP �9�}����f������u#I<�	��g@gdt�gH�ONO�;i"�M�B44�E�*��q�[YXH����f �<?*8_���0~���-@>
g�)R=��:���}(���	 -k��'b(W�P��WӨ3�ݘ��*bO�O�]�J���U3~�@åm>�����i)��.x$}մ79�x,��b�|G\m~���=D��y��UW ��1�����3̑���(���S�L�����
�R��QK�p���G%.:�5��	������B[��̤*�w���[��u<?��1�Vc��1��';�K�4B��YLYÑ��7���p�Fr,�]�	���[+��*0��ԫ��頼BH�z�쨪+pS�)���O��Jz�s!̓}He@�TTUA��޷��b�8/��w���p�MN )7��(���b��xu���zg�:��[�]��b;��E�#����遡�����m:Z���xǌ;Wj�T�s�g_�"!Y�����	�p[�Nގ��e�<�Z���kk���\ ��њ,�H`i��E;+��*...MƍZ��sl2n�'��~}?[G�;�G�Ri�?ފ;�*0s���������<%��,W��4�Y�Z�-x<�ŵl� �UmwrF����2ט�{���y�20PH3YJ��d��)9��7�B""�>�W�,à�>�?-4�+��d���W�>��x�.��u�W�Ѳɮ`��fc��4j�����%�4�;����N���(��Fff
\��&h�&����*@~�T���h'�%����o�bl�2dݩB�y?���͚Jd������&�8��s���^eR��j~��Ū�*V�Ek4��2��٣�`����,PV1. (��k���R�����Fp��ڿ.3�$Au�]�iK�<���w�<,A��U���Q��"����_�����5@R�p�3A��z�a.B�x�ݹ:'G�x}�a��mzͺ�F�ko����Q���M?��@�%����N���d a�j'�pIL�w��B�H=a�X5i�'}��`L��w�h����5�t=6�z��{��B��+1aS��
2������ō�n�~���|ౖ��F�A��]��{1)�}�+y��55jyyy h�V@���{�����WPw��a�Ǻ�g�������v�,�	8�
I�ɊYh�v�{��~�8�\�
��$�PS�Q����{�@��W�޾y�������5"2�2���xu�����(p[�� *u>�|ՖHiT#ΙcC�FE8H�a�����d2fj)N��ܸ���V�;S����%%_��X�A���:�]S��@3ն�����0�ɓ����C�5Pj���ސ���w�sܣ֥���-�_]7M^��z�3�R���ۙ3�-��]�ܪ�A-��L6���מl���+� W��ӫ:��#��><�@�"�����w�eM�fLh��5�� 4�/	5�]����$�W���d!_889}����奤�@ǣE�=;^ǜĸ�9Rj�_��:�?�9	ss�h;�Zb��]�}[����G���������i�{C*P�����2�MK0-���Gg���ʦG�}Y	�0���[�j��ϔw�T��0i�S]̤��(� ����m��b�5?/`�M��98�'�-��3w4��G��, s�mK;;�<Woӕ	��7y"��Gם.G����ʒu��PZ�%�(�7�fD:ChK�0�����������Q�nګ!����߿���Y2���剛ן�m &&4Hح�E����#�*d�qQ��f�Sv�@2f���RN���A:��Z��˩xy5��.�M��XQ\6��P��Oh���{�����q��+�s���v�v�J�͠{���q�"��J0� $����9::����i��fP���D���dZ���Z���z��#�ZE���U��+d{���b-�r�0�C�1����r�>K�{�P/Z��Z��� �N�L[
���+��ؙ��j܄�1bz}yy�W�nw"�:o���o�#_�*a�<mM,v��@*�@���[�gK�K��T�`7�Rj!ϖ̯���Ԓ��e�����ި���L3=}�a�#�t��Q�Rg����5�U{����MH-�ġ�okEn���&X�%�e!�������ْ�ВF�2�Qt�Q�	�"D��)��hB^�t�3ri>�G0�dXx���>/E��[��/���!�#bI����**�+��\�D5e��d����،��b��I�Y��2�kU+`-�rO��W:9����k3���Y_�u�zWY�XW�SD��;�{�x2%����V^q�r�7��#�(pqp2�r�q���J��,���-@����AsQ��-�fލݽ�,���os=�"��H�ϰoEv����xS:�ϴu���N��Z�#�s�	]��OQڀ���"Q�-�c�I�ÓӺ0w����o@
-$:�/����g@�����]��?�����T�}[�[b���ʶXy���F`Y1K*f2O�E?{���?%�g�BXׂ���%���h������v��q�r�>�TC�W����z���Ԁ���JM�:0s�d��f�n`�s�ׄT�d�LLֆQ��1,��h0���ɕ��N�����8�� ��7Z8��͑IC�n4d�����ȗd	:�|�C7�,q�g�Tp8e����"  @CC���]�g�.cl�H�$��p1�<�m�Ɋo��W��Y;���P&m�[��><���.��:#E�U#^��H�k��-�'� ��b��VO�Ji�Ւ/-��r��l�:l8���f��iV�o!*þL{\\���-(�.����a����Q��ꥆ��%�=L74� ��q$��
~�t�y��蹜蟂�1�9�����T�SU?�W4k��%"4?�4O�.0�+3��c����~���i��&�l��i�P^.~G���!��~0��Dfo�7�'WUqd�^%�׿7�E���
���A�g��֣*A�%����h:��^�Z��0J�uI�!j̬<\�Ack�U˚�et��z蓌1b�EP S<��z(��X:���r"h��ړG���r�����j�V�wxH���[���xw�v���D����V| R<�`K�4��^^\�� \5i'��-�׽��3��vE��t�d���dε
>I���+<N���k�Y4����VH�E�O�c�!����Zr�{��RM��h]vvv��"���D��+(D�h�}t��ԣ��� ��hn�����Փ\]���sJCMF{R�KWƣ�vFp/8>T{\ٻ�<h˜o���%P��:z͚x�%�r��=�v�N����H6?�a ����4e~:T�? [}j��pّb�����}�O����e�*���n��7��?y{��hX���i[�YmYʕ�*�2-�''!x�z����vo�֞�sqY�$I�$�?���YZL�RTi��׏��~̤�qB�����n�����$Y���uԋ�m�F㎖��{�*��ü�	L��*�?+� 77w�w"],����,@�g:^M��R�������|0W�F��t���Y��*�%#��#."St�ۃ������:S��K���\8�����5�������k��67<g��pm:�rǓ��Z8::��o�X�h �h��T��T���ռP���c�ex�}_������H�����wnh]]��� -���P%DOO_d�*��BD��X�� P`>�|��� �=��B���wFaZ��n����_�Z#S��J�_��ț��5������{���خ��f�^^^4tt��=iO���3:���D	�j

�fgiU�zu�4j��2* �8~t��"A��L��Zہ�����~�l��K\�V( ��i�b�}��c���`Fȅ��R��q��G��v�f��og�/B�Y�Ӿ�w���\e��F���`V���Ȓ����s�[\J�im��b�(���礥�SPP���������@7� ui:J��/egW��f]ee�ȏ3f�`��n�������Y[Q�ӝ"-� Vm���`r��<�˥u�PhvN�M�퇙YY��l:��bҗ,�a�?�DU��L�ǟ	�T~� �5O�T��n� �)��:�w=��٭`����֥�-b�l�|�}��)quyaa_++���U,h|�o_�v ��&��40<|���/��)sh�z�����E�?M���Cj7G�Q��ja[��ܙ�^ǏH����ŝ�p{��tS�hqq����?0ǝ�@���e#a��%6�|u1˫$�n���k+B������DO���q}��x�uK�4��6"�ێ�Pו�c�>~�<>� �?ߙ ���ܿ�	�ד��5kS�J���rҢ�������Y�^���;�E�2�'���֭����Q�q5���/�v�`wy��ĄX#���/���2�����2�V)Ě���/����¤�:_��#^�7Ş�6+����:�g���ǆ5_��z��"HX�i�|O�����n\�_Y�}��g�f^�-��B1�7���v�%��H7��|r�yLY����&_7��l��}v�*,���#K{�WZZjğJ�s% e��ֳ�d��w�7�����7��YlO�e��X"��E�䭭.�eg����	X>��n�Ꞅ�ǧ���~�ғ922��ݞ�g~��ʐz�?��Y�#CI�X��1��������p��&���׀>{_m"Q����^�-(f��	L+�v�7�J�}!ȼFFF���+��]����	������4?WII��y�3�rw�Y�ةli��LDO/鼿e��""��z��ٞ���r���� FB�$��n{6>�=t�r��ü����L�8ρ���Cۋ�	g-
m�r�Ȃ��$ ݄C�.�{q~��@�4:�a�DbX�,������C�	���IÅ:>f5��>�פ���a{�^t��r$�	�7�o��E��	�.˯�����p9��>��,X���$|W!_-�hT��oSi-���˿s
���3�烼F�+�b�˫�j!�>�-�HY�WU&?~�|��Z.�Kc�,��>��pXH��������24�F��X�RI�sI<�U��Ŝ��B}�:�����\{��j1p�W��4(���&����uj��͔�� 5����Y�E�&�4{:�pҹ^�Eȥ�)(�OY�_��Ž45�����o�r��B�v��a������!�u��1[M���:����?�q�=�Ӭ���uc)�##"��!�� ��A2'� �~��rJJ���xtJ�ޙ���0O�=j��%���f%)x'!�u�U礁R��j��Gm�(�(f��5�4+a9�o!�CM�B�����{�G�(��k�����9 R%M޿O��w1����[[[%�K2��Ur��nt@@V�D-{���ή�r�q7S�� �[F��ƻ�1j�Fook���LJK�l��Y8(^�-�������d��fN�ن��YT����"vA���q�n��v�/��q���cP��\HI!s9,#*�QMmX9�յ�L-�6Z�{���,����'@��տ���)GR41�)(�[��ܑ&�ֹA8 �I����`����e3e]���R��v'*Ǥ��$����R�
m�;���```@�P����/���%��t�õ�J�B������C�
mN�R?��q(��G�pyih�8P�_ժ��S.d���8-y	va=jC�cBӄ�S e�����S�А7�;p��&" ۃ����w�p:W����3���I���8�c��hH�������Ud��w4�o
��v������yA^�}�Uo��>8:9A���/��	c[�ݟ�%	�j%��z@^qs��*���Bӑ�_"6u��� �j���V	��p�J�`�E x�c����������5?\Ǎ����3L�Ra˟��m���\B�מ��� bW)�����"��$j�9��C�����Ы�������tUʳ���F�
���TJ�?sV���TJ�Q�%�`�U����� �wJ9ͺ��4��
d��L �p,=�V�'�$P�p��"�@��HK�u��܃��0>�O$��bqz��W-j��)����{��t�t�_��YG9�՝�����/r�I98T�/M5z��(7U-T�1�>(6!ДDp���Ǫ˷���Eڵ�3�P�A��c��?݆���iYHH_zS7.�rK����c+F'%o����\{����vM*��m'�6�+3?~�Ḵ��|�.�G�1���-7x As���l�^��]Q����;h�-�Ɖk= ��`�L�o�--�UK���Pr�fWw=����5�gU�=�4��#��f��p��r����Q6jI�����!݊~颢�ۇ�	OH�S�h_���N�r�I@j0R��?ȧ�w��/I�x6ٮ����-��g�ߦ�@��1I6��*���,oo:�ܺyq4)�Ҹ�� �:@��L]�z�X{0�/�r�bL ]��'~�� ��5fS�[B�x��t��`KZ�l�el����I4�S���(Y���[���*BB-��B�B�	U�9h��������7���8�I~d���15Ed��jh$�Vl���Ffȏk�yE��[��3��(7�tx��Δ��	1$gv�ڻ��� a645�wq����-�[�P�l�u\���y)��؛�p�ފ�n�d���0(�v��	*��X/ I�j`8 ���Ը�yÀ�𸱻��UP 	�Uf����o�R">��Йgna!'3SH@@`˞#�ĺ/]<lr}h�ɧ�n��F��8��qzW͢������^E�6Ə������bl����M����Ms�7`Y���/��!hg�S*|[m�nˁ!���D�[ng�DF*��+-i��e���y�p�e�8��k=���5K����P����(6����Ձ[�@��2�$��O` �0්���~���4,XT�m:����@�cc\Fn��
�I�g���MC}��5�飴�:���;48�����ᷫ����{0�{$�B������	�xIl-~��Ƃ��	<���hg5����j�U�M�I��瀯mE�綷�w�����A�U��v��9Z���]^]�377��~|_
<�� ��̟�x;��w2T����SV�Цk��H�:�o���y��-ؑg���ْF�ϓ�����=�Z��jU�E���qza@�C�sP�bh��<�9G!/������|�ɒI��>��R|a�/�ƿeI��$���(y?V�� �ѝ���3���P	��#III���sVByQQ(l?.H�x���4���8B~@�x&���'�Y��<��)g6�bJ���3����]�����l���޽���-""x��v}"π�&
���i� 1R*���#5�x5�?t��b�p��<��MIh�t���n&%���Nh�kpp���k /XY 5䰘r��eβO��xps��l.{�^M��l�* a��� ����؆�`*	�6���]�����»)��I��hwe���0��a�N] ��`*�Enx~v�Rn��tq�kZܧO7q���Y}��9�B�- %����
'��"hց����kPA׬�9 ���{��GG%n箦�u�@�Ά���-���g@��K/gl�Cgl%FaW=�Re�\���q��[��)�|�Ғ7�Mn?Lk6[W]ҫb�iW��; �H$n����7����&=׹#������)���AR�J�RQ�d`UO��r��$�|v�V�o�l4a7܇YoL�i��첮��e�������t� (R������<����h�	���}��%�����N$B��'�ru��L~�q�~�W����^M�g-�H���p�32:
0����X��l;Ɏ��6��V�䝡��\����0�a���y���
*%�����J��I:�
듅 �T��`�ѳ~'Gǝi�GP��g=$�iDq��d>�����I@�w%��Ot��H�8r��<�ċ_e���p�g��̨�u��on�y�L�=mA{]���8�bG|e0o��b�[B�,_�O 1��6��i	uA==��溔):k� �AG_��w��v�e���fgcc�Й0R�Vӣ��#:8��Uez{ߡxЉW�á2�V�w��%ҢU���|ȡ`))z>]�p��G�g}��nb$�{��3�.,X�6:xN��$f�i�xe���]�n,����͖G��P�l��zuQ�:25�R��)�����Eg�����`����������X���ǽ4�^1�1d�z�L��,������+��f�#�0�2S`{jZZ����(�-���3�r<��_��"r�邱n�S�5E9�Őw��K�"I@.J� ��bj+Sp/��:04Tъ��ϰ�72*D���2kW�'�ګ4�zy���V/��ٹ�^ׯ� 409�軄���mO��E=G,.vC�j41K\�2b��+������>���T���P}���%Q,Y
b�R��Ԕ�����cPSȶdX��c�o�Ru3�b?άB��'UIߥ��p�w�˶F�}!�2^>\�Eh����Y9�<	 _������ͣc��BN/>��سW17�����srrv��pȘ�+���)&<z���c��6n����
�����QXA`@A`W	i�	EB�;T�:TXBPR�s�!D��a:��� ~�g�����}�=�\+��k�G@�Y���u��Nn9�]s�yGA�2�vonA���|��rF(���}�!��'l�rm�B&��+f�2 E�{q��&��ۋ~Mj�o˺?WX�@7��q3��V�� ����������Vj���@��
b�c��+<@-�m�Ėp�N4H�y*T�.d|6���
V:���nn+_H�\��q���\*;�E�C��w���?5c*���� ��ǧM+|@@ �/y-���M�Ha��"�;��	;�v��o� bf3�!�/�v
�liyB+�k�cU � %�4��q�S������5$$$;�#���k����?䈖|	��q��y���Þ T�7�	���r[��$lb�S6��5�.y�t��1���D �M����9tV��osW�w�.w.{=�(٢�_��@k�[�B���q*��x|tJMC���Bm���ZF�V��#�k	2�3����XĹ/He�t�(9C~Z��i>����� ���x����� �iB�e��$�����\�q���+��sN���{?�%+��)�_b�ٸkW���j:/�+(��!K�ń>�=��%6��0���a��&��~��Ϝڿ�� � ��۫����'��?� 1Z�*���I
?�؏��(ԭ�.�p	~~��z8���S�:�Uq]���^���G��+�S��ώ��&�WhY��=~��rs)�����u��hu�+�s-`'�.h"�%��W�T
��E�F�N��OGЉB��I��$e��П�$��dU��ma�%���@��͸�{M2��CPm�[M��){g�h�i��W��Q��@�:.qtT��TL���=vJ�_)�k.w/#d�s��Ma?	b�Y�dr`|�-��%q@�@9��kf�h����o�=�g:\�Z����Q����]ETW=ڔ����㺘%%��珃]o���|�<+/�����eQz��㛞~�ƃH�˵��<�Q	�ѷ�Ԟ9�-�U�='&��9� |�@՟ W����p�E�=�vhv�Tj,�ݏ�'dA���A_�S�c��Rt���g�UH�I��e�fݔ�h4�ȿ��@"
�B�+1��_�I],Fh�bq����
������zßI�HC�!��.ۋ�c��\��YH�ɵ�R� �#n������[���&C;�����mAپ#1��ֲ�k@fj+ЍѤ\�c3�V  Y�5��;���;� %�\~e�U�[�x��Y	(�����}y{�ѫ���n�[��9� R�l��FF�ம�a%F�z��3���sF�<׫,���
�(����+-��/Ҏ�|�/Kc_ov;��ڛpӧ��|`��h3E#^�ͤ��\��_��m��azt���.]2���t缴�mj��x^��QHL��(}q�UD��x�ɳe��(�yG�޾��N���_!���$0 nO~��ް.U���� m��/]��q���Ȭ����Xf�X�,�Zl�[		�\����>��S��Ijkkc����N%��������K{�(i�2_��x��ˮ���Ίt��u���|Hq,M�.Ӛ�9������� *xK䤜S�)Ub7V���a3�D�A��X����˨ͫ׷��ѝQ�ݓ���J@6�AOx&˿�#Mf�9!��yu��-��E󮯭�9��(����~	6\�k�'ٗ"� ���fs��V�8�t����l������<ɻ�CVj%SXQQQ3����|'�ml5<t�_��N|��YZO���������-��kЊtY��jeffR���\�J�h�W��̭K_`�\m���Ye�� �0 X���h��B�~�����\�r*�W�QW�܎'I����}��m���'�vdm�f(����J� lY ���j4�k���Bh��\�|>F�K���v�*��W�Dڗ`��5W�{�����ņ�"�����;{{qU�_����W��h��+3E���%tW�Tb1���k��#������_.���A~�����z}��io�y]N�OV2z+V�%�M�,�9�sM���A 
�� 	�~�֠8�6---N��Vkv�X�p	�s�K��U�$��⻯�6�.e N�����"%%-��.����T������\vz�!� h�Qh{��k�ϵ�˲y���� ��jۜ����u�������*�""����Ȏo^,8!��1r����5W��U�6 [Z��������Kz6QB6n+ ��#��ҫ6w(_��G���t5�7X-_��PWW7K�N;Z�&��>�>�\ᙙC�M��p��D�����-��i:�}�����k׮up_+2D�,?����c��D�hlUdd���Oz���*�@��U-�A}�SL�/$�멧�G�&���J9��ը�����mY��|e��쬠�b�< _�F����o�g����7���'�m���҅�O27�j�xԩ��>�U�X 6g��U���t=�-' P��ҫ:��.�~���U�΢,��������..���{��/���N�^�_@ @������<|iܘ�s����0�TĀ3̎��/�|�{-��w�Հ���XŚ��ug��nL0�j�/:���h|7"���ٝ�:θ������T؛.a7|��*�^jD��of"{�h��O����VV� �궯A��?������3Dw��(�R񸸸䥧��8��kP�?�7C=9����~
��: �u���|�-��}�A�e�!�<��0�� ����:Sⵉے�r�ܧ.����rv����{�����sN���[�l�G�tc��c����'��
Pe�jM<�ʣ��R�i��6]�}h�"m��T1
m�d�;�������L����}���tͫ)��.=�~2���) �k���Jn=�/(�K	-���o�Tf5��,�S&��a|~˻�B�7%C�4Í�P.5p��&$�g��UX}||��
�Dv.���C��===�8e�J)�P������f��Ѥ�b�ԍ
�q��_D��əW��m�����ӥ`������,3�'�Xb��9K\�I�����M=�A^����}�<�c��� �C�\zE�����Xj����=|����?K��
C�B�/��3Z����x�V� �%�����h�P5���ik�4+�2@@-��X��;!l�#���#?~���h�?`YF�����L��xN/Z.j�[�W��rF�ŭ�|nx�^R:m�,�U:s��̘�Xx=�����Gx�w�������u���bK=���/�m�T��8NC57����1>ᮁ��eu��\���>���>�ap�tw܁�,Tx|�\�¾}u��P��u444������`D[��;��t��C�;k��Ĭ�i.ĥ��-���@��l����g��Қv�#a�%~P��}%��>�NQ���o�'�O�p}mL�̶ۘ*r������u���PϬ��$��mƞ��� co__AnnЯp~(��{�6ŏ�Z܁�(e�$c��g���;p����b�0��@ 	խ�g]N%����i-[K��ד{ע��Mx��mu1��]���"+�"��O��:�<V��"�R%��yg�EJyUs���yd�t�ߜ��x�ĺ	q���kM�L4��[�STȳ{Z2����Rq�&+Az��������e�~.{��� �t?��ث������]o�
��,�Ғ�D�/@�b�W�ӟ��l��~E�C5[��c,�������F����ކ��������{�m��
x��M��e�k][�Y
L��rG�����w�~�1�X���8���<�~�XSǍQ4-�BlO���N�!H<�f7n2��X>1!�+����C��	�6���������* �%�iR� ���xyy��=(?j|���.�N9��g)��bn��?�A�dr�M|��n$�8� ¡��Zx�[Zק���]����C=�Xm@�L�
�g��t!�J��e�_���y���3I�� #,�
@@-3�����Q�ە9���bb���,�5�i���M28/���Tm�=通����&��<��pjq1��H�J��UXZʝ�����p���~s@3E:w���n\��C�߽3�Ϡ�D�vܾ�C�x���A!�ӆ��Dy��Z���l������l�ΝV��;`9Y{V�D��
�	�FZ��yb�h�{��4�(���M�~�����)@ 䓓��ի�� ��6M����	���O����j�?~|

���
 rc3��S r�B���1%h��{{�r��>���z����F2�w튑��@��$�|�q�������4&�SC�V��l�p<��ؾ��Rf|�Z���9�eu�b���d�~y���P��`�A3ʹч� �M+b ������D��y��U�ۏ���koEў��Be�y1�����=�Z���@���(�GXT�ֻ<_�K���$����S�
��b}����P������)���N�f{�s��
����6�-�V�	�{�`R�X�3���Կ*��s��i�'�r�T�a���W�u��j����s��RTVnn�H׸���s�j?����tܦˤ�'��9Щ3�.iz�ȓ���R��K��W�=���t�;r�A�΀�؜��5yd��w���9e�'�$��,�������r���ӭX'�T6����W�K�~�մ⹁)��m�MFG���"�{	�c��!��/�	����|�_�,lY�u�Pf�+j+E��ת�G؍il2YGCmB&6I��뉩1 ��f�bs�G2�	��Ƭ�E����TU<���^ ��kL[��w�CO�<	hȮ�r����p��@%��5$����Pg&�R�R��Ï�L5pGM�>X\Q�l��cW�k~���9�-Z.{xd�"�|��
L�`� JB�E755�ހ�nUp�s��D�L��I��zL�h�q�~ )���E�?@��	�
�ק�0���/0����Ⱦ��a���\S��Ʉщ��Z_�|�R��^�g+���a���o����mf���q\�Ts����������t|Fcͪ�55��FC���G�Xo��(yJ �1���IɃɳ��~'a���������	��p�M�r�` ��E�T%������,�gE'ם����
�@�p}ڴ����g��-��d:|m�'{	F⟧�jj��vZ���45}D���2y*��G*N��HFF�Y�%�d0҂���ϗ��m�lVE6�I��<���A���#����~LC��ag ?�mG3@̳����7cK����&�J�G!Ղ6�RdVJ�͟��-�7F�,��J���r��ϊ���������\���4��K���Ю>>���;+�V=)��B�bC$�0
�������)`�Y[���T�*b~;�;�ד*����o�#��A jU��˿�h��E`c�y��݃����\���rp(Yu��3�{�4�@� ���o�P߹S7��~?:��v98��"�������;	h��?�ʎ�؛= ɺ���i?���:�S�V�_�����b���\MP�X�ho���	��ӜS�� ����wG0r�sPx��~J�����+i�Ny�C������A�{��6���m�@WAe��So�n]#d�P�Kp�t6zx��>��R���J�y��H,�{Ǟ�d&�9�Q��hM|[�p�ЧBwsZha*�mmm����r���R#.v�sѧ��T�0�� ��ŮM�e��Z���]�J�~NuI��������&'��O�]#�b���eu�GZ���K/� ���f.��چ1�V�t��%�����#�q���>.����#i�V� R�K�~zP�t�Bsj���Qs�ՙ�D����gb�zz+-	q t8��<c������%당����_�jr7�O��
�ܘ��m6�t���0�"�� �g4�!DeƉo���u�������%��m�;�iil�>^`ޚ_��C�0IZ�u!��ֶ��6�뾚�.��U�k�BJq�	�,	�����>jض�F� �Mջ,�SMZ��K"ƃ?��U�"Ϊ���f=�Feo�]� o�T,ܱ����8�|�|�s�s �l�nE�;���=��-㍫P�����4}���V����!�N�ZG�CϪ�)��q�A=tWo����0)5F�j��^�k�/�N��A��6|y?�}��.���]3g+��I!��G� ���d߄��& 2�d�/���}���3<5�Nq�=Q%Xw7�8�ٛ�w�և���O��6�
��04���oBB��	hiE:��_Q��ʑ�W�Dj&=�W�%���q�2���ߡD�9G!9�2B7�D1#EW(���~�� #2T�o�	܅�
���M9��!򖆏���I@^�S�ݏJ�Ee��M2��7DT��A3���հ���P�/q �`�����to�\7���:r�aKDUom-�tM��rk�̖��:L%����
 ���'��'rF��/���u��Gwɤ�]7l���zyii��A:& �ol|\^ ���}[������/��PNz�'�<@	�p��/���]�:C	p �c��GCn6����~�v���xI//��|e9`��A�P�j�q�Q�R� �����%6�s��gz���\>�txP>'��	D�4yy���cW`*���ꛞ�w.�oI��TP�=���h��Z�D�tYHA �J���*_��Y����#j��'M�->c����m���V�����G��H��Zh5ED
z��м��˽����e�e��ֻ�%�$�2����2W��&3J�CɇP�E2Z�,��TBR��uIWO��S<�������ff���wP+���ܷ��&�����s�,�����2y��w-�x���W� �]�q߆���jƋ�5y#;����o��X�_&$$,����0��o��jV�ag��@��5�[�
��><q�D6"5�$S[ .�ᭂz&�T��o'l3~���$���R.�����XĽ	�T(S�?�j���'��!"��>����~���:9�'��о�u~�*��[������]k0➜��{B���
9J�"ǫ�����Z�����.�w��+j?0�ΰ��o�@P��|VΠ)��p�ky���r��wtxSխWW��]���X���r�mm	@�QA)��Gc�J�#W{���~ǸC��&��'n�8�����U�8����-�"r-�{��׾��&��៖�gҬ���r�nvY�����';h�=�GYZ��Ą5�D��$ "	Ll�J�����E�
b\^�:�n:������Q��笢���=��N�i��33��z�>�ی,����,)w���2Be���;�_���@�^s]���dӿ��W�t	or�%��C=�(���q[��蟩p�o�C�lBb���Xf�%(*(@�����m)	h2� Iy������l+�"�گj.O���ꏡ��S��/<�S^ {�l�U�p��i9�^;a�#����I�����*���F	 -��1���;y�c�Q- zɧU2|�5�1����� X�&%%]��G�-{������m4]!����R2<�_���dQ/-�$	����+ ����:89�ػ��� ���ɛUu��h���2ޛ)x�7��4v�C��������!�?ۡ��3��v+���\wu@��N7"V�|��Q(�u\OR�t�IB��Yf��0�"��?��$P `�Ag�7Jo����I(���B��V/�	%����>R����E�6Q?#n��T)�o����|��1Ҷ(��6���*�sobW	�c�*�^�ܣ�3���e�<'p���aM?����bW^l���#���3�S�7�{M�ԏ��݉~{U�Pϕ�V��n�0G�ޞ��C০�{����:���5�`�K�Fj�>�])�n5��p8��/������%6�* -w֣���,DS�x�+.�G��E�w M�W��e�MJ��Q���.�(�E��w��ם��!�����-�����	hy���l�;n'�_`nN��ןN�6(���GD�<�K("j�_ ����W�;�ƅ���7�|u��u�5W*d�VπTw-1&S�p5�P���ӣ�Z%0�>e֓�?���ho]�+ ���/��AOJJJd� v�8�D�JN+��[Xu����9[U7'�g�.��&܀'�h(��_��|r�б8m'p�T��=s��,=/�M�<>@m,i9e-�l�F��ĥj�`���Z�;�]���dVc�L	��W���H���C�\��˳�#'��s��y=�+zQ�zg��\�/	�f�s!�}8�o���Z�Ǧ��<]�u7S�s_��'���O.���եde̬sv��eX?��/OZ[閨�ϴUWd��8SD����(�Y9W�ڡ�h�����
�8�\s��Qy�����dd^^�pZX�hyOr2m�.n��}�Qv{�Y�X�ʆ	��o���h�r��:����_%hԕ*On:�X��I��^���+B���8�Z߂��ƴ�J΂�u&aq��s�!��z�(���^���4����\:P�R���W>��y�/��6j�ebbR>�f��Ps~�Tj9�~5��(:�N�����ӡ菟b?~�Z޼��D�Ip��bi�N�"$��߼�l�s[h����>������TP���[�b�4]���X̄�ƠG��vla_զ��y߇�'4.E���?���m��.��ژ����*�z�N�(�����c&Q�l��9�:Z��&KT~T��1�u�f��|c���P
�-�������+�=vJ��c,���dTT���	<�cy�W�R^���yj�0^b&¥3դ���\��p�YpEPh�q�6�NQz���*���&�#>11{xV�CQQ�������On��#,L��������"���´���|[r)���������=Wk��s�|�䭭�X��Ӡ��96ぶ�4���~���s����)���1t����Q�t袰�>>��呷�/�/{>�B���s\8��gs؏gR�3m7,�)�F�\��?���i=�5X� �3� ���Ne:
�/�m�Th�4���fN�	����E �/h�nz�{^�7��߿_?�!<����ޥ<j�}����NY�'C��������<Z7��>A��yz+D]����9
������";B�~M�Q>�G-�5��R"��W��7AǦ!����<��}�,��g|��'|�V3���o�i��n_o$~��5��"����ji�ٸI7g���_� W3�`~ۙ��?��B/���Y ��a|�XW�݊T�3��<C@�R�s+mGyD�V+���s��;'#�����{��/����˨F�\RRצv��h�Ǿf�--,�`n�`fR3>�2����A�+47*���՗��Y�L���j�N�,���{A\/������b��}��Z
�&�u�� �ֵ�����1G*)+#���L��X����}<�Urn�͈p�pu,�sy�VXdW�L�p���&�����t/Ĉ<��!�W�41��h�z�tX����	i'i&R��Y����h�>O$n��)ؕ��[3�jg!*��د�/�@�w�G���7�.8���	'U��ї�46��7K~�[��.����ؐeP�f���	����(U׬;����潴����}����4�'<%ic����/R|��K�[�/��2�4�%������t�?�-���֠v��2��ٵ��Ղ�C�yg����Y6l�#خP>��yT���V4�k�y�4g&$5G1��ѷ����d�E��a:� ��?�Xo.�8���9�M�z�D���e��NP�Q���W(�0'>.��į�SJ揮/=91�/tO�E���#GU�J'� zk�A�}�߸|?jz�����z�1GFFf`ż�{��i\��R��Pl:=@D�����k���/�~5u�N����V�T�;���4�=�/?�3>�.Xj4~�ߌ�"�L����	#v�a,zsb}���9���Q�e�JE-���1����u�|_��3�֠����������	�6�$�?I���]��+���|��u{8�����K�T_�(�fM��ҋ2'�d-l*����Χ��WJ���ti���1�<����(jV[G7��m�t����o�(�<��9ڵ�nh�ʏNAn=��ޕA^�Dlu��"�i��F��j�~�3��|ւhKu���(Y	:os�3�5���\؂�$mr~��I��u~N)�ҳ�I=�Z�O�7�R��I)��/���b	�+�M�����xѫ�X�,?����ou���LB��Y ��ݳ<f�8y����L�*�	a�fqY��fh��kUII�'Cǃos���?X��{�"r���\�e��	�sݴ�ŏ[�d2,R<�O�MҒ�������t2F%{'�����Y5Y^\|p��7u�3�鿯rw�� �)�����.�?���,�����DD_�����CR��E��b�w��ق�eZ����Q�Yff&tpxtT�q#�Y�
�M�����s���<�{]�)H�hyK�[=���6�]����y�lyg>��:�|-.<C�%,����t����^��E�I�R���49�,�xd�bO_Bo�e�@Y�@�;J���}^��@�J�i1��^_,F�i���Z�i_c`�Q�`��i�(��參@\k���QZ֩���Li��]�{dx���<ϔ?�%�ޘ�������9�Gd��	b�e�A�s�{���(�NN��{y�(�a~nnGu�g�J�P�����[�)�߆��U����3/MӒ����C�yQ���)0���I�b\˶�*:����KxXB�a%�BJ��NS��V��} �R��j78�(4��`Ek�0���Q��l���{E,�Xv�v�9����[	����u����:~����-�e��V� �5�9G!��:�R�o��l�_OT�:��+����Է?a0�
��b�`���
a�������:�b`Cd�A�L'LQ�E��	9���+Dr��=��[&Vv(i�2�a��rL��6�I�v�}*����V�s���h�S�W��q.�	9
�!�iH�u�wƵ@S6���G"C��#H'�G�U�9\�Z*D�`�:ۯ�z �M��ٝ{�K��RXZ��UzkQt���X�����,�|���K�[��N���cKt���Y��
L��R��A�uO{�k�ʁ����d:O
�9^g��6����0~�}�I��$�����Q��5OvBGQ(I��""'7W�\vF.����xſ��ۡ���&�`��~���~K����?��3�IN^,u�Dz,0��2(�ĩ.if�=��e��F�?.���J:���o��BTkP��}#�lOLa�w�����p�<�	��31''���gW�>��9�4l�6W�PX��_�et�)T]�?.%'P~z�cdd$ݾw��y�s�+��n��6�����Q�9hP3���� �����J��D{ �s�;�A�K���Ax�Ό����{Ή����Z4NCV_귨�%����	���xG[FC�-�����6������"� ��	&�������������U��!��qv~��b�#z�l�����p�n�,;�߹ j40���c�70X}�E��T��vy��+q�t|0��L |�W�/t�� �ݴ�D�20���t��þþ��F������0�#�r��;��F�&��'�����^�]�a��U�H cGb�_�R��]5u��w����#�宓��f�C�|���/��s;�;#���L/?��G������`�/	��8�x�V��%� ���mv~x=�C�$��4bh�b$~�ޜ&Ee��`*���9�B�:�9�^{ˋ��e��V	��&�\(��k�"u'���u~F����꿚/��Ө4w��]�rV����JB��j]F!�����;VW�T݁Հ��!#d���?�����ӢGK�x��l�x�FX�<��i�3�#�yx2pZ�y���P�*p>�w�N5�z>�%CM��GGu���Z���
ݍ}y*��i&*Fw2(�[ֵ95翉{4��\w�w�牊3��z*��ӄ��۔!�$���fuN����ca����lJ����C��+������C�"č*}�Ӏ����������uq��)m�a��/�jg���j]� _����dq;��B�D����J�ˑ�]K�]� ��Bi�D�.�;�����vK��7���>=§��Qc�^�i( 3���5>��1!��m���׏��KU^)B�y�
A�\���.�Q�+���F˳������,Ӏ�`��ո�/_�Q
�J�~�\����Q��]|<`ݯ�a6���3��G��~�$ϔ'_���u	:)�^�Y��x��We<뮾��jE{��>�.���K���5R�Ni�����d/uz�7�=M�'0j6��oE��փ�f�r�؟?K!��`�~�m	OB�N6��/����=���Lu	&�Sz��w	�M�Y+sQ���Q7�b���)��x�$%��<���V\r��po`غ\]���bk�ͱ�Զv6�{�X�ɹF��k��4��t!#�tlw{�enș'/M��JH&@��%o�|�9�1�
�Ha�m򡦦.X�[��8Cgĸ��;�G����4ΘMIB�+��jօ�������te�"�� �ʔj����s e��5C���~�����9h5�x�M�F���>!7T�^��/&�N�e��$�|�q+,��?p8<�__��p�/4Iȁ�82e" �c_����@Y��t@p�$ә2�, ���N�J��YXU�|�4|���B��BÑ�����PV��tr�����,�
�9Q�lY�õ	�6��)���B'f�$�_Pa�4����f��ù�oX�h��[��v��]B�JP� ��"�*CθX}�ꃗ��o��w���٨�^g��B"�6T�;��t>5_���r	 wyΘǿ��%&"0�@�c
k���쫸\~	�<�0���a�'���3����_i�N���o��g�X4(��+�!�YM8���`ζZ?��'YEst���ѕ���9���+�ش��P!���6���EF���H���~M��*�p8tt|��@��^�wh"���tJop�*YN)���4oF��ΰM-���O3�`kF}9B-L:���'BX�5�S2i���}�\L�ŵ���6�2Gկ��}�J��^p�P�A��Q��`�{���*W�v	|��F$v���Ȧ��^���f_��VBk�T-��h�Vq[�0������ ����[z#c@�G�ǽ���d<Vˏ���۷���]G�0�D��*ӎ�/O����:�=sa����%u��(����~:���p�x�
���**�!�
�m��d[��[����'@x�>vW!"���
_�GF;�њ�6��>;w��kw6BP����M^��bXM�p���f��I{8K�KƹW�	9��GvP"`W5��p�p��y�M���+\@=�>a�6����.}�eX���%ӭ���Ac-����/�qo}[�̸�&\zV�Re���f%�k@����^p����E�7��2�M�}�)/B������w��{�>�ӓTh�=�mR��nge&������o������!@��pu'�|�-�w�r"�,6�
���^��{��	{ƨ�/�?[W�*W�*��(�P�:d��?!�� U�p�?��3?*A#$������������5���㓅Z�����]�=l4~�ݔ�/���⮮���ץ��SL��Д����	��<\���%���4Ȩ��`�/v�U��\����~�0���������S���4���W g���eW���G�W���+7ズn.������<�į��-*��rg<_:�:;�L@�����9�`������U:�u�L~�u*N���������x�Q�ή��#^��u}}QΜ�+|��z M�u]w)����9^�� �hɂF
u�G�|||��YlH��P��&֚qßU�UW$���u�=�3�1��h�R����@\{��gʾv��.���D��V���B��W�Q�S]@򟟐�J�G�<��&���6��Fю6 sU� ͣ<�3a�a+ U�E�̴^%%'G��w�h�Y�R�&&&���P� ˂�&���L�uN%�ӳa	��=�=l"^[2�ΣD,ഏ�Kh0��z*.#������DН���8D�Vsue�b���meC<zn��������B }?74�7Л�J}L���1B��H��8tw��o`�V@�����WBэ֛P���v�\�84���#ګ,��*���8R�O�9�{�;P��{��Sl��q���v×�5e#_�(/,"ҭ�fn.��>~� "=�(���X�:5�����4 �)Ӵ�����H��w��nŋ���dʙ��}�E��Jko��Zr	��$ ��Bm�����e��NC.���v��I���ț������W2|��n�,��������%�UPm�< ��K���r�j���[�Yʏ ] �vwיv��,���I���I�i�O�|�j<��^1�Ku�A��.s7�̌�q��$&nT��8R��b9 �	�:;%�vQ��i�o�T#�9
Z!Ǵ�ܲ>��%έ�o<;�����f�8iy�W���ᖂ���T�T�f��+Q�U*�����t�:@�#���W!�Ζ���X;��-����:��hHd���k�3��S��N�ﴂ��*�ȿl
�Z�r�G;����q3��������������o��v>Eu�x7ǚe��}m)��E3�9Ң��ͯ�Q������ps��?6�>PfVJ�������X3nO*а�r�CM�5�zB$,tsk&��'��8����G8���*uh�_ٺ�&����}�6m|�Y߃*tQ�{�Nrv�"�3�!%#���)�I����6�.�,Q�&^�-������̙��Xe���lk��==k	))#����K���m�SD�q���՞omgg�k�No�:�@�˂%e}��->|	��i_Ӎ�С��6��H��о�|$�8M\MA[����x��G��@��E}T�-�Nq �w�3F���<K������)1^��A5='~dA���2o��&��ع$is��<|F$911a��k�B��c�T����!�JHDD��0����d�z�/>��%���$F�k؀�� �+?x�m��ۂ�x}��{�tW���j�C�Ru��/��?�!������x�B@� �����mZF��j�&���S5j�X"����Hڻ�^6Ϻ�������$g����at�i��}�UTF�(� �@��`��]�q;U����B��{�����i����ǖ���{�Q_̣x�߬��>e�*'���΁�ׯ�?���fK�ק�
���GE[f����$������J@'#t��OKLhDj�Ԙ��XxS�ax'R����Bw ��w5hF��=&��ݬ !	��5er�	�H���>�H�2��\�\��	,Oη�9ǁ�+��~�8�DT�T����]N��p�+d-z���P��)�;�GNNN>�4�];�c7��O�������6B�B�|���Ϝ?�bl��L���g֏��R���^9M��Q��I�uKV�o�+	�2����u�����E�U�udј\yg=�Z�k�l���pS����[�l��,��i���_�������Ϙ	Q��
�����<��|�4�S�׏.q/.-��a�I��5�R^�09�	

rX����mf��=����-6.~��:[�GM��n�.dV:���談6^(_�A�7w؛��7��%��V~�P�э|��a\2��M�M�v-�WՖS;{�GM�-	U��0�Ǐ�S��n޼	��kr��>���ܕ�o�����|��nC����q^-�x��?�F B�-��ݰ�.�,dH�+J!-#C�r0鵞o�)R.ho��1��(Ǚ�D��	q���s7/�=X�pf���Y�CE��g_�n������j"w	f�-��|r���,�}wL��O�6.Tn"�|�J��ի��_��Lk/
nŽ�����ucœ���xz� ��tu ��|{5��],���[�SL�Q�,��R��*�z�m���w�E����m
9������O�H@5���� ��&
�K��eX9_� �-
$t�I����]Y��5�MP�
�E=��{�n�8��Y�C�^���ww�e4��bz�'��%�+�`ħv<)���eW����=�g��ym�>)��$����faa�{����Z{���p����.���/vTX�* �m�����ָ�\�M��>'�eJz::y��@�Px���/.��$�>���t1%��k�9X�J�H�Z?�+��^9�{� Z.F�J1^юS�V�������?br��3���b����ZՇX]�GF�BG�᫈Ɗ�e�v=����9S^U��G	�D����1������f$.�L�G��,]LO__n�]&����\,\p0[KYc�����;�k�a�U��egg2[)����w4BK[Z��x�:�\�ة�_9�V&�Wz�� �?e#�ۼ�W�}���dffV�Y�A���1�$�eg ����s������;䷉�)�2>�O������L	)�We��ލ_�~o}z9K*5�2����>%f{���Û�C��C�:�89t�99i�x�j|Β+��
 &��^��s|T�7�sX��ܷtt�䫕,W�,����) l�t�X&S��:f�������>����{3v�5�:* �l; �y�) S�����$ԃ���2�����u����T�j\Y�r>�n8���N`��Gj�K��v����~#?~|R˿u⬣ma�p���8��!�4F' �n��}�T�1.�L+��o�aWLED����Ǯځ�		I�zh������+b��{/b'ȚڟK+�:\�Pܐ߃�B�c\��K�Q0�~�(��a�5f[�IG��2"��knm4�l�K�5&�b_kO���j�ʁGӊzj\@\b�������8B-�����~0����sg�pZ��_߰���IM�
�m��v���"\d��!��2�*Bv����lb'��4���0�[�z�/m���]�q��|S ����MB<�m���+<�w�������ٶ�`��n u��l��ӿ ��!7��q#`�ç-��w��;�g�G'��B�V>ՠ
ɯ]����rB�33�Q�!�]��7���-�{{	).�^ϙ��{�o�q <� �İiC��|��<h�~q��)��]��lx�?���Y��2sD��A�e�Zy4Q��@D�R:���d�z-r��|��̎ҟ:U�(�}��<�>vs3M�p�#/��sKˎ]=�b�2�a�����V������gcu��zU�fvĝ�!��� ��k��Ŝ	���_2�X��[oF�4��e���W�{�5��ƨ�?2���7��dY��K�\�U�?	��WW+�=ob�4�M�� ���N�i�e�g�#��z�U�D�%�2dXO��l4�pl7qSP��j����֭�o�p�R���zR6f_l �ӫ����� ���pO��]�T��8��#�"��j�q�'G�f��+8�u�ʘ�ړF��0aaaK^�J�d��TSid�p���޾���SzZ�M�$�j8����Hz�b�+Ā�x����k�����hxbb��.j5��Ғ�SU�UĿ��`X5��oߤjL �U�}����N�$d��u�aMfM;ꂫ���"��T�w\Q@zG�J/�C��"������^B���C@D�I	�tBB����~�%?�}w�9���}�s��H�UKo&�e�Ϟl�}���l& $T����e�TY��������9�Qd�̯�GTp����(C�\:���Qz�q��\�cy���ّ;����ؼ�����%��	:,|��'��CoK�)��pD�j|�#J���jq�:���[gQ�_\RRQ\www�&����2~E��^]`��!i�����2Gޓ�f���$�g啕�_�̅�ea�����a���_ �XI��]�u.�^V��[�o�QÄn"�I�}��N�1�� 7�Ã��l����nTʲ1�%�j���Y$0z��_#\�cC#��H���eM(M�0����zJX5�w��s�'L��ҏ����4�D0���p�Q��@l'	H���R�ԢJ��o��q�0*+ݒ2�!i�$ͼ���t���/D �Rew�.�+�>(�����'��t?;���\�����E��z��bf�߹�08j3v����� �CxWb\gIH%�{y��N�XD�o_�~�<}�9�{������kc�9p ��N�$�J�sC �4;;`��,��q&{����z�<]䔑����;�����t�E�Y���P�SE��ڽ�ܞƋ���,��O��ݝj%�j��:C 5��p���7�VҠ�L�a�&&S����j�T'n͜{�\�����hZHXg~f��hg{{�����I�f۠^��h�-��`I�LC�s�� n-d߄��T���]pdI�|\��N�&/`���_~<���~o[��ۊ
>|�sV�E�w�τ�uL�?}M�Do��:���D�9�������ꇠ���I�����|
�K`2{��N!�@����;�T:��..�����Md��y"�G>跷�2�ʋ�+볲��%j����c(�1W9���>���������p�����vN��Q�h�����67���0���Oa|#Y߆XܥV�3�4wE?��;�QMoo��^G�pIn�_�*X��;T� ��A7����
� �C��"���3g/.�d�Ũ�� �87��ep�b�&���r�^����/kNtWF������rkRcufZ��c}���[�+�g;⅄�r �Vxs�Hw��P�\7q�o#�jܳ3�V4�F��6sA)��bêvA�*�b#�&V�����e�D�4�"}Sά�_4:F۴s�j�d[ĝ/������>4My}wf���9��4��Ѩ�����c߾D}����xM����Pa��-at@�gyJ�\8G߂��1�o:�v������u��|��/Guս�S�$�aĒ���b��B�ޞ�~�p��p�J���;]]]�׽K�|fq�~�b�Ĭ�D�N=y�~R@��{
�H)%%��� �wG ky�HɌ�õg+9�"?߮�ʂ�˘:DY��#�a*O�Id|v�Ī�q>r�U^�Y}zNEU� /O��<Z����k��p�L*_܇�![�����i�I 	�a�gΎ��4�0 A֛�Q�WI�-qƾ�&��w!�8����5~D�4�*[�NS�)r����z�Ɗm��g�aLӑ4\��;���N+s�� f&&'������G�^jz�.+����mY.dGgu���!��Ë��o@�r���Yn�^�}��_�v��U��$K:C<��nZ7�ҴP�g����\�Ipț����-$h������� ZS�W��oit6�9��4���;X�N��ϷsrR�R�])���\M��a,��c�eQ��9pt��p�k&%w��yڽ��謫���ۜ	5eX�߄cll�r���AqBJ� ԥ$��*D#��?�u	@�(c�I�J��e�����S��q�5�{B	-EA���'��G�l�O�=mH��U��G�K>���a��@`u~�n����\-�k{�o[�4;��fu=?k����l'|7T���Π�����Tϟ�f7���2n��˵0kkP�'��2���&�`��uP|�Sv�a�`��]�3u,�ք�@��\�� ��2t�w-l�lncn���d��4?p�Ls�C��s�!YK�ok�WC~���Csq���g������`f�郌4ws��EX'»L��ߒV�n�C�)XE(�)����e��nU<����n���ɯ�$�-���UiUQ&h@�o<�B�eEmzU��JRB���`	7�N�_;Xa��8˲�#�1X�]��LP��z�/���e�r�I:��Xݗ�qPe(+y5j��-q��]���Ď�Y�d�G���
��56M��}�g�pU��B1t��&M���O��t��e��/0X��\�:�!�"&,-(�8g�j�V '?�u;�����+�1�݁������i(��w��V���u�G�,�+�#������Α��ϑtk���j�)))��46F�cu�ɇ^��݅��1_=�������5_)��p�]���7`���V.���dv�޷�P�(]�}J���IIZ����i6a��. �����*�������a �����������%��ס|,��ϖ�ĄI��������e�>��	�i����ЪR���4|�h��
�ņ�}/�z��@�P���4����!�Xd1`Кyʩ���pY,!h$�����A�w��Vby'�U����g�{L.y�����H"4�%�����ydVV�����-�<��:C(bG,�ߣt��4$R�jj��C�(��Ih*�Χ�����\��bKb;��B\o����q����8�$�p�Mi�Aԋ�Bac=Ϋ9}6�m�7���["��2c�.\\\#�pC"E�6�=)���~����+p��kY�����<��@V���["�uj���R�V̉�x���+.4�vd�-���5��L=n^"B����GFB�� ڌ��54�T����<"�`����⧅z����?��W�SN�<i����Q�xr�D���>E�Gj:��Q��l��ɭ~-�rhI��L����N;�A�ѳ��8}������h�{u�gaN���A`ͳ�J��ޗ�TƵh��i��X�(�#�s�E�-CwP_u\�1�YTz�Mq<����/��n���>A��p̈́�;�++g;�(w��Gி��ϧ}����Bj�Wb�3w�}Ԡ�Y6!����mK��
���1�(:�3��J�b���t��b���3��XIUG�������~lnV���`�wQ�B�if]�h�~/���D�i̴��f��>�Ӌ�`˄
�|Sw2V�����x�Ӗ�F	]}iV�ۿ�X]xS�g/�<˚��nM�
3Bl�`�w	����
5Y}�h�sX��8@��P=��׍�v@ެ	�8,i߾�H�=^s;%����k
�}�Tu!\jw��%���0��u�]g�d���	`9W�w5�NzgQE���Ź�$C���N7��rz�BmH��q'zdS[��i�
����q''i�G9�����<��ı�\.eN�r��X�W�V�.i|Em�#���c�ӵ9��^��)�)��[��V�� �rP*�Ø� _����"��^���lo8(���K�����6�f������/�2|���D~��>�Xw�/�8üߟe�p���=�*�%(-�����궐 �V�,��bF��`�GDK�ߧ�jN�����>��l���åB���1�u���6�6!/ �_�gB	�\�3����źBbbP.?`ٌ Tmh�d�"z�F�3����ln�i����o2��'l����߯=&�ӧ������2(��.
}%L�<��u�a7�n���y��ꆧ$b#X�
�ߚ����<���([�<�+�s�������s��_�h�Tt�D�K����*���*���@�	�6���R���k��O�D����C���J��l��:<\�\e3ۑe�AX��Zf
��93sss�q0N����"�	Y�U����7��i�W)�������0Tj�D  py~�#����G<�ħ��e7�m��{k-�|2l�,�`�Y۴�zTqLk�p�G(�$���4n��3(w�E�5�}��ٚ���q	����MC�0F��Z�ow��A�۴@3��QZ��	d�=�FE]z���v�=w�� �رmB�Y9y���P=_&�j�P�������*s��W%S��R���uwG[�}5J���� �ѣ4� ��v8��� ɺ����\d����Uw����GeJ� �(h����TNS��R��%��Z����A14<�J�ރ�K�>��vZ7�S�}im�g���o�ӣoxE�z(/Dz��#���ɸ�������Z�J���?v"j��(��,�*�<�τ�R�7I�v�1�>:BͩJy�m�.�vԿp��[%���AC�Ž�4=@��_w���X��W�$��ckҀg��c����ts�?�RT�q�lT~?��p*=���w	�x��R�s������e�U'�@�]ϴ��$�"��[#���w^��<�ӀQ*��bXz}��ߍR�⢢��W�N�Q+�b���q`8�}�p.����[" �(��f4L}��\�]��U���M"8 �w��m�֥�:^��k�F7�)�+m�ėo���Ti7K�*2A������~�#9996$�ٿ~��'�P[�s+��;1OS��ۃ[S���f�R���(�����| a���]p0��^�Sк��!���4�cM�Z��Kn����F�x�+�a_��IM������\�?#c��#++�_f�vE�����:���x��ZE��.��J�b��DSW	@영��w�Y�S�u��Dg��r2m��au��������Ss�l����͜��,�М|?��QSV��	G�e��[.��J�+ԓ����A��}1�Y25\�+VxS�07���a)\d\���Y"��.g,T�ݔ ͍�YY\D֙���ct����v��^��x
�,�#���xϱs�OO@����ۖ[��{�5�-;G�����E�i��G�#[�  ���y+�Ń[h ����6glE����z,��N�_%��������퇁>u���-z/3��sgEչ-FC|�eУ�U�顱��@KA��g{ٹHs�t���Q8��61t�6ko$�rZ�3� j\�g�V�Xa�$��@����w��t�w�UǊ�����Tˍ*� D ��}s�]w��r�G�F��Y$�*����0#w4XL���D��.�X_��3�j.��d�lE�{����f�O��hll����-pf�:��H.�fl5��8U�����,sG?N۠fɃ
�(�����ClGױ$�^x���؏-���;���f?��g-�OKJ�r���nm��H���i�[ڜ�vV��ꜱ�2B��F}0޾)����ǁ>I����|��r��ˋ��%N�ܥ��|����VP��1Jl���V2�-� #޵,M��օsk��$��1�)��r*],!������	ɳ��Ϝ9s�2hVF�D�ߑ~Pp��Xe�i��]�ez� ͓�^���xs���� ���pW󕖖�D�KNA�;������g¶���%^�&�?��M������w7E���\��  +ц>*b,"�#��\��Ãj�3�Y��c[.�b�b��?��������v�wĪJ�&K�j��F�'�$��TJf�6���c=��&�kO�.������#�<�Ӛ��������+��n�����.'��O\�������muDĈ���!�5�R q�D"�
}�[�`�~F:Hm��Q��T󶠧�Q�,����WF��c*J\�ۈRk�b��z� #�5��YjM�̃�ڞ������4����I�X7ť�$[l[qҞ����cb�*V��\UĔ/��u���RQ�'�eE�}�����˥�q�Ôp�l���&��G�V�ǲ�v��_|�˭��>5����ig�i��r���@A��6��	*N�k�+O��t��%5k�Pv:���"17..�m��H>��-,���M������9�?��/�병:���e�,�Q	]�I��k'*�,������"�1��/K��	+xLɄ�� �7����m�W��8���^�mm|���������x��P��q��� ]��|iU.���?3����=QNb��&U��H���6�J�Ӂ�3F���xxx;E&��bw�:o�#I��'�o/|�0}�/����NC`��nٛ�D����\�LǸ����'
�1[obTbq�;�{[���΍b����x!\ _�hl�tE�h��:��ٌ�<��P����7�gM�@�2�S�p�Umŉ�]$"�^��ޜ�����l@&+**�	vn�����饥�h6s��~}���?z"�b�4��2{12�7/�|������E�3�=ҳ���B��a�i���w,�(-��7�/����L�`�kz�{x��##KvZ���da鋬<<t�>���ަן��h�.-@�:�~*�ʺ�o}�D����*�rz�k�}{�y��S�*b�"��HU��I��W���I�*��K�p�ƀ	���n���_hg J�仨I�}*�#�����4ռض�m���⼴����
��ws�r��5��d2�� �۬�?�c�ҕ.��L�X�)I��&�:>^��&��}+j�vd�L����Alŭܖc=NWFO�#;��	 r�q+k�0�^E���2��G��񟐜�����X���l�;��κ�4������W�|��'����lB�#���.��1-wH�Mէo�˄<Ѐ�N��!`�W��NU�m���%�F/[&�BA���m��Qk Y�>�彄���HV���k��(+`��-��3"�������`K]P$��Ь����D�ؑ��10���iZ��j�">@L�&�J.�����C#��{����;��ڼ|�yP*���{����"�	��%�Xׇ�!�e��)���k����*���أm�~��������V��D��Ϭ�N5C��wv��3L1K�_��x�{UW��S�ȸg ������5�?��ɘ����#��\�z��-�I����=�@jA�����É%;L�������)UI1|K�����}�9C`�~&%(�0�.�
�ٚd�ܚ�)Y
T��~��0�"^a�>�XŜ��@�%�>Q"�J�B��DL��ԙF����|$���P�Z@���76������)��N��&��	n�Q~*��￙�j�����|�)�Չ^i����:3YenJ��twFv��8C������r�`���`#A�u��#��/��J6��A==!A�l�Cx-���\�i�[0� ֥�hv�j�'��x��ㅟj�>�9�rb#�&'���Kd���K�=��O%[�A�Е6�5V�͡&��Z4$�i�ո�l�ގ�+W��-\sDq�}�u�p�0��V	�co�Yvs��m��5�%ٸ���I��0r�D�?�����b�9���Y�� ��bccC�u�w�˷�������TF2��1m����B����ݐ��{4�ׅ��">�H��p��N{{{붡ܯa"�L%⬼��k�J,����~�1$����^Q���WӏQ?Oq��n1��'IڷI��o��v{ۧ>�h����鵒ޠ'��E+A�#}$���o�����߈����:}pC�}ˉKVە��9-�裴9�'}�1	>?l��V��H�YHٰ��1�S@`fo�}�pQ\|<�䀔�hl�TxE��;}x(;�B�O$��L�%�?6�P__Lʓvbz~���H��	��0�%�j�.���`��7��G���1�|�����"��$���)����1�b��������9�s	�o
�
��k��?�Eyy�!��J�|���ٟEl�r^����x�sd,�n�(ieeu��;s��yI�T�⦪��>�۾5q����j�$����_)�R��bMդ�>�\��;��9^N�Dz�2;�[�:~:��}�����&  ��|6j��{�5|��>�dlYq�4���_%�Oݕ�Bg�o��́�S`�<K�D�m̻O}����jxX_�36�.��o��q>1)�=yO�S{��4��I��SZ�*��)@)wJ�rfOn]�;�g������)ԁ�q<���@K�$~�O���?M���|D�0R>�!?5	��Q�%j����Zg��{��<�\�[P#jq�-amN���U���56�?%F5/}�( l�я=����D��	���`o{n_��0J�s�|熹�IZZZ��,J1'3�b"�������� Q��r��g�K�Q�~�RLO�TW��)K�z��&\��@o\����U9�|6�+�V����ݲ��d` ̊�(< w�D�W��t�G��]Z#
#���ЃT�w��_i����Q��Lz~<���J�=ҵP��'�����/_H� �]�7Tj���2V�S��L���s��a|Y�ֳ���VhL�uZ�B}���s����&{�#�^��D��`�5E��\����Tsyx�M�.I�|1�s��G�*R�ȸ�bWlm��������&�j�z���44\ש
�q���,@����ј���VsW3��V�ޭ&W/�X?5��0���,%&��(���w�h���)�M}S��|���;0�C룚��p���ٰ�����{����K�+�z6.g_	�HJ�N��)sL�0��~�8������=�O��i�,�?���988趷n���AxD���|����j�������ǎsչ�|�)$��B}{Y�dK����6'|�a��(��b���	j'�a�;U���ջL'z��M�yRP�+�l��Q���$�S��lu�vP��r?�G��#v(�},ܡ5�9��O�U��MA�
#Jg�b7��Q~I�`���IHe�TS^>�Į.����ܽ�c8����nc�@<��L��ڇ])�Yx֟ߴ��V�W�\s�+J�:b��vq`�d-���
�_{��rt,pK��jqq147Rq3k�ZS��$cAN|#���~�|C���#f��n��/����SE������VHI����/�2X�菝%{t�Z��L�1c���4�_��vF��i\�s�����E��Y�͐����
���\xډh/�$K�U���iERu���S�9�o�J����vNjy}Е���\��ܐ�"h��$�yuQ&����6�1w�j|���>�i���2L��7t����^2��5X��i�k���<]��E<��$^�,���Dj��o�d��?�Xt�����%������[�$�t�X^^�]�����:�{P���(�N��>��#j#��I����V��G�½��e�Bd3 N�=΋8�p�j��z��Q��iaa�;�ș�L��}?���4��T֯s��t'�A.�k��������҇��p�=D&'2�����Ya(��S��b=������F�7���o�KF�M {{^�	��)����y�t��g���{Wk�>.��@,<�l��Z �4��f�*X�&�P�9������4�C��z��\}�wNT�S��<L9N���
����ӡ�I��y�Ax��újb���.�E��J�}q��e3fek<+�{-#:��H{yq@����Vyћ���KK�A���`�6��',��� o��G�KXGlw\Y��4�7���yw����% ̎ﰀ���|MJ�}����\�H�؟Y����l���I��a�栺c��J¯^��g�|���h���L��p,�S�v{���q�ē7hA��
<lm�R�H��wa}�c�l�b��VAn^��+�}��Տ�qk�;��V��X�
`D����:���������BrVS#��;B�L�i�  �9(�:��Gl1����T������;(h�f�����	I
�u�����}�m�~~=؃t�:O��i��&��&�bkq�D����hԪ�˟�.�%�����8֪W�s��A��+T�K᥅�[���FY ��w�F�k቎C�o�IL��U ~"��S�D��wu����T�ء�^��1W@��#3�]$9�T��s�1F䇸���m���.��F���.\w��P�������1`�L��t��'��"k*m���pY�ć8�����U��0��6��=�;�]]]���$3��i)�����y�8��=vdh�q	��xI�cG�&/E�E@^������t���0;�r_1Ҧ�	�Q���ϟ/ǲ�&IL��oM�{
��L��u�7���:�+�[(���ZE��DE�W4�(��'�5�{w��}����`���:�A�`M�΢��>@U�W�G7��"�3�0|\�e	Px���gk6��5���`I+�2�~Ocg�M1+����EW���E �����ee��4���,�c�AAA��j�ƈ{��i�$O����|(�y�n�bbZz��B��Yk���{�e�w�������<ǓJK^�VK&�`�1�S�|{�Y2�Y�(�c��mV��4@p<?�֖�B�F%����cv_�!�iLP����W���$ɂ-|gML���J8T/N],�M�d7�975t��|W�<AqP�d�����,f{�n�Ch�=�W�_	�[#�^�����x��ڀ�;K&�І��胣mj�!qw����'~�dwc�7z�A��ބ��t?��	�M����@��T���y�M�����FZ����i,�����(�p �����
�`�C��'�_|(X-���uh,��Z'�?�ځ�L~t�W��o����P���)�qO��I+�(�ơ���֥�ܒ���~�����lУ�����V��+�ż�8����	2q�)�Ѣt.eQ��#gqq�y��Kz�Y�= �P�6�-��5�x��OPk�����R�>�?�X �ޚ3����*�I��h\ N��Y�������ej,UY��Ej̆�aް�?tZn��k�^����{~�Z�$�P	�'���}�f15`�j�ܯ6�!wI�,L����&ͭE@H��=B�g��3�w���[�ߏ\���I��M6
����{�H�}ë,��r
	�:�m����% �Vi�\��1m� 饤���"��1�r ��y��Y��QFzlll�VD1M��\?zT�K�������H���)���iʈ�(;h `�Pҋ���
ƹywd$Q����mO̗N�z�y�u��2�V�x��?�\��m�����װ�s��Idq��;�X�֩8+>0�u��uը��Y1����p�U���-��
�C�8��j*�j�<#��V.���_���A��i����p��~��LC��6 0O}Y��z�}*/	s�4���;�q��I�wj,�4�g7��#I[��~�4�p�c2U�������g:7hH���c��<��׭5J�:��܎�}�}k�B4�Z��N��CXX�=�8�0w=1��P:MP���Ly$Ǖ�_H�v�at��g3�|3B3}� 3nu�v����ş�n���c�����z�e�6|�E���:��q�i�������I�=�ܳ�M�?L�ݥ�4�nB����������ا�O�_4�M#כ_?���tni�I����LȄ^Y�����3s�	$�;�����̮���m9c�^}�+�����!��̏%!�`����c�@��iٷD_�k^c&l�������P�i����*`2{���!%Em���Ƿ�K��S��UO�?��^�";�����H��AB�ev� "Cw:���\���q��<�_hq���C<9o�oU�0�W/Mq���>�HϏ����B�8Xǲ๗���cθ��2���߷�Ӑ�8 ����;�.\�RVQ(r��y��-HpW#U=8�N��a�W͛�Rw,�_��NM��`��@.�����<�SK����7a���BW�l3bM]P� ��ʇ����H*�9:+��j�nma�������ќ#9�a#e���V!�HVh ��l�)��I�u�<3�h�欞��Z"�rGxz���zM��}��e�w��Ɏj��qq[����D�C�2�� CuO�Yw��=�;}�T�R��fT'M�7r0�ڍ"p��^+�O����܊�� ��ݐ1>�z=R �?�K�����(9��������~�=�� ���Z��Z58|)1ދ=�:֝�N3�y��D9B�h���K�6t��ebT�?Mw,�l��JH?ށJV�q�^g_¾
_�QW%ïW9A_�=��9���Gr��⏜ZB�q���9�)�t�q�F���:�z��]d�� _f<���xd�L���>9��a�Dg�u����9��CVV���
v���i��X���SfC��U��a�q��Q��vp'q{�\�%����`�Զkm�`�����V������,bGY+?�-Z)3�3�^�(�
To}�W���No�x-=�x! ����|P̓ӄ�H̍n����;�`����:R��9��=e՗�o��q2�܅��𧱛e�	:J{���+�Q�z�i�)G���!���Tx���v8h$;����_�ulz#m���`|v�M�B�v�d�_��w��f3�P>ii[�1�M��'���.<R,�����;8���H%�v��<���Je&��1;��Q0r@��eH��T�sZ�-0��s
��v�r�fOʾ'��C#�ʭ�Gj�$�(s@u�~KZi.��e܅�^!�f�,�W)fV�c�V���:\�a�	A�+j��G}/0��m���x���u�,���`��J�4����c�������=m���
سV�S����=�\N(M~Rom�4Ec{h �`��x��"�6�Ǥ��	v����z0O�Ȇ>xꑦ`�
wb����]�A�w"�}q���[����f:�O�o/��3>�;'G�<�ä��z�T��5��h��L���I���e�e��>�����}�����di����2�w~��/ѰA6��~�����]�!S� �������&�q��ٓ��	B5�_[[�c��N�DPa�)Mǳ�v�Q&���D�_Fp��i��$SRR)��b�yz4�J��J�(��@�f�*C���D��6w�;\{{�Q�zV���(pG!x�d��E��o�4m����>�}B�1�=<16�.�Df���#&���vRVd��h?��b{��Q*��n����C����¡��������[��N˝a�h�T6��/"5���5
�geE
������ж���~~���&*J��~W+�Ϳ��$��KѰJ�l�����9��$��ZwBr��<�����HZ�s0�G$ �p9��#"�?��� ���&+��Hl�c��G��b
±��b��Ɛ������� k�4t�����Sw�i|G�um�W-15�S��G��Bܜ
Ǵ���	�j�X���,�r��j���� �*�@���jCi���n@uo�v��"���~\	�ng߶���B�ڈs-`U��oa�18?9�܏9�W���̱�;� o����[���n�B�nV]MM����^��l�����klJ��i���3�h7��n��3��Ʒ"#��r�2еUw���z��Sl���}�'�(�<�d�j��3�{NV�p�hhdȳx=���>��zr�R������VHM&`ݣ�N�Ed�?� ��&ѥf��2,7���]U������b��	���T�%�]̷_ɕ�;�?-C6�f����u��WV�9���؜�1�{7Xk�*>,�~Q���$aq�j�\�Z���:��s��)�����X~ԯD)�k�	�-V �r�T{�4t��C��%H@X8�M������"~Qz�'C�����S�I��e��|�=�_��޶NCy�FA�b�r˗>O�e��,z�D?Eף��'L�6��C����ق��$OҐ�!V���m.��@w�G�~���B�C\��C�#,�@�LPZ����0�v�T���R�P�PճR숵�raf���{�5�e�m�u���,��`x�]�P�A�i��E5��4,ߟ	(Wq�J/=��~4m]�U.J�1�+���g.�.���**M0Z�u>�s�$՜{���v��Q|�S#��پ$L�V��"��*�q��4�c^(��~' �N��#��8�*`
���<6�|���p��n�+��7`v�>4���0����Ό��d2��lÜ1�y3{��Wc ���O����JG7��/���ן֝�BbG��a-/ŝ>��gl8��'u�N	4����~��YGYA���WQ	���H�����'��?�C�9���M�ָ+����r�,Y�n��'s�,c���;���Ii����P�R��������$/��N�>��Þ��h��b�\Jܸ>�l�?S���(hl{U�qR:$���ׄ�����/ߟ��]~.�o�u�Y��"�#m4��ۿ�JJ[�nG�;���^�HC��u��~E���?�?2��,G�$i��bnͳ²31���s1]��<��hV'Ʃٴ�1�l͙bH�;j��t���B�m�_���Z�q�O��1�����;׌9!I���Z�"%4��M�Q���m.K��>?UvJkm����9�#v�agc��[�IWCC�k[�޳z���[>���1#��xƥ�Z�2w��J�kb�Vv;����.��rxD�l��`��ዚ1�\�3OA�ZZZ���<�I�=�Ex6;%� ��娞�h�8[��+��%�
�����;s;��|n>Y�� *�VMu֚��p��8ދ_�I�7�!{ qw0���SڥN_s�I��;�����阎��w��i��g.*"ۮ����]ŏ��Ȭ,Y˺�]rv�AlU��������w	�o�d��׉*:��bM��ݡ��k<�A��U���e�j,�z�t�3M&�����Z���ߋT�N�ɲ�b��W$�RW�%?��ԼH@���|�A�Gh���py���������D
��]"˫�ulZr+���H�s�T��1�ϥ8OrM�7��%�'�5:���^�R�!�@�����{f��2�����£b��Q�2�ؙ$ҽx���g��)^�ڷ�oy-���+����Í��}�ظ��2����$9yx�cBk�p<=����m2�zp��Q4�
��}�ݲ}�Mv��o��$��;H�޺����i�W��S�����T��_���ꣁĝ���`yi�f��cONs�����Q��snL/����ͫǟ<�Os� r i���훂�������4j�e;�U���tл���ɋ�#h.�Nc���:��"�axdda]��:���n���4�uZ�V��8�"o���$4�䓡���r��KI�x��_|�{��8�aw͔S�%u����S@��@yh��a�}�?��܆�z�F������;g�8�;�b�5�� ��psn<���Yr4;�U
ܑ���g{��Wq�֨�����)_|Gl9j�FǷ�K�+�]~�|[�L��p�ߴ��ڲ(�������}��.���ut؟z�!�I��-A�	�9ո\�碣]���Y[snyYJ�<����W�a;�*��\�@/��Ų$����yO��@�O��hh��Ԍ.�<x�=���@����I�Ʌ�P��4�i����/�?�; �of/�~����³���xGkg<<#b���caa![�bE�˫�vw�hM�Լ�s���ҡ����-���R�q�C��1�3k2��@,��� ڪ�2s�=L�5�\������s��(�D�	��n��W��]��n�r#E�M}���7��ݢgԌ��:��
E)�����ɦ@���j�������Uꂀ�*,q����2S|�>y1,��Z��S�F�S"�c�4?t�\(����s�%|�S���o��e�9{Ѽ� �^�y���˧��n$(/m.�As�S}Hb~�}iq�,u��������V6Z��ܳ�k�xf�mK��aWeh�����wu�wR�If��P�Y�Y����0h\����Qw�$*���)ҰA�]c�0��%��"#��F�k�8?8%�����3�����d=����j$ԔʥRO_?A\Bb`` �Er������f&_)�L!�=��hydYHn���~�M����L�ؠ,�H%����t`�?Xb�Uu��� �ao���*��;`K�!҅�g�2��'s�sVK�r�dC[�!���V� ں�V�Z�K�H]VV����2n�K�ݵi�H|G���4[�ᶻ���oc#���>52�51GOE�kfh���2G����޿�l^u�6�ר�����I���Z��ighJ輻�5�M�;���:�Ö�g�C�vt���GJ�l�� NN�(�<��+Iv;[oΏT`������ʢ�Q5����؞d�[-9.6�\�Q���Zφ�<��������}A�����=�B?R
V]��5 � � ._U��fݧ?v�)�뀫�bԝ�216�y��A�5��ţU*$n�gn�`�����իW��� �L�R]s������4��S������^�e�z��PC���?��x��Ĭ�W�����@֧t��d��������!]	7ln�`>{vhE&r����\�c��'��8�"���xp����&$FF���K��=Е���lii�T�*��H1z��D"ָ��F�:�QW����iȹ��GETz$�X.t�l�Տ�;>�g��+��{[�m��2��A�ZZ1}G@�e���YL�p\�* �H����׿U�1��\�^���*��׏*ZV+k��/^�---}�"`���kL�4[:M��QƝ7}�����َx5����<'R���r$'���Gs����L���Օ���L�S�!S���v�_�C����ٽ���k��me����6NN�GGGׯ����y{{;���;���$��±�[�� ��a#���J��o�Xo@��Wz��**7�o��~*(,tݏL阅���>5�,f��#!���߱(��\6�"��J�3נ֦�;�X���Q.������hGG'''�S|�#"�/��P�-��h����j�c�S#��6'I��"���Յ��KE�Y��E�#]���3ϻ\u蛡� ��F���G�����������9����@��N{�Lm#���5O�_M���ڊ���o�z+��y|�<e���G,,����n\��zf������T{�6��� �o�����j��*oP�f��N�3��LÚlG'p=11���1�=��W�͙�4�a��Q.���_����P0z�{O�'f\_����
��:���\aG��K�+V6�8/�����;/}��S��N�ٙ��?X{�e���,t�g�{��"�M3 +�TT3w�S�B��-K4�@��Tn���o.�Z��	 Y]��,�I�טE\�������w�xoWd�5���s���㯞�����7Z��"�>��jGˠ~�u0Ah�k�<|�^.T}&�99O���틞���bb+c����G7�O�%^I������@A?
�/����L���7�$Q�GhM�Bگ9F�]��PhVͻ}��i
���m���1;~�������6�c����:N�=�Ј��� *
J�����}o�EU���JǉTp&��ǘ�0X#<)�}�d D:�x~��u��	 ������T[ϼ������6�BXR�;N�${�ul5�2����<���Y5Z�����Lb߉%�9ɩ�I�n7k�j����sI�+����'}�BDi�q����� �z���aRBZJD�D@Z��F)�Mw���l����DE@$6!nR�- �����|��k�sTp3�ֽ�{�̚ƽΩ6���
Q���v������Y`4������`�}h8�vw˵���y�b�����!�A��d�d�IQΝ�w�W��<�QG�rEp-ź�eIA�w�����Q���%��-����E��v2��;)��@h����/��%jY6Z�X�SW����Z��#GI���	��k��Q�v�9j��z���w�T?�W���qE٧�W�VW�n�@�F��<�)�(EI.b�S��f�A���k%[�"T����u��	������C�\�5�P��,!
�$����ö�|&���R�>��m�E�+�&S�ʕ��ҷۘ�	�2�<�dx��gp�R��oVW_�a(�a�䗾>6^��y��D!|�!�]��iC�'��f�5U
�6X��좏����Rj�q3s�����;Wάx�%Oj�2x�S�M6��������K1ҟ�73�j� �[�'�����tM�"*TZv�K� �m 8���\R����5j�(r���A.��MjР�eM_w�v�*y�p�\��"c���M�5�����g��+,++S�=�O�S�1��T��d��]Ac9Ӏ)d99�_>݋ �d��$�0GX|J�%��f�kuI�R���s��op�ۼ�6�֝�1��Kb��갦553����˪�U+���ګ];��hZA�����^(K ��r���E���2����X�^k�}��WcQ;�)w=�P�:��J�!�u�3�fNR��.�vnߍ��}Ĩ��#^��=����Էc.�!��X���)�و�n����u��+vŬ�hڝ�R3$��G��Yӥ��6�����Ư�����g��v��8͊��Zo?�a��*D
�B�+�*T�z�EĲc;�R^n?U�`͔�h��@�kG�$q�ɓ��N ��K�@��Y��<��@��ڐ��-�I�a�r����s�s"��[�a��Z���;�T����+���gR˭,F9�w��x�~r˃Y�t�pB���l����~�:��p��/K���*�=G�vM���D�][L���r@tf��y��%I1R����`!�7���֗0o������T J�{v� dle '��kl\.O�k�E5[�t ��ۨ�ˉ��z��>(�>���ш�����������&�TT���*��Z[���d5??�$��t�p!��epӊ:�/�ֱCb���[���[ќ������r����Yf��g�~'��ss��*O  -�0�:+�<��Z��^�oOOr|���z��;0%�m�����|��T���ד�/���d`�`�|gyhUQ��AHD�
����{_X��<����|��M�i��Hz1@0'���I��~���-6����0(�:����ݲf�1��'`�x_�3�%#��D 3%����ˬaي�~�i���F@m%ɎC�;R���p^�Z�!@{g�)Lbq��)�J����c�R "�s�V��C��0Ϫ�m	b�/�@�@�@�Y��n@P5�.��cT� l'�>�4�k��'�W]�v�(���C�uT�j���h�ܱ���ぐ���S�����!�:W��������Ӡۻ�V	;��I?;����5��~q�J��"S��~󴰑�A����P�~E�����o4P| ��=��m�N�ΐ�q��=8�V�S��k��ؿ�зl���v*�j5n�#T�ǩBW��Řg�Vpp`m{���k�'��ME�}��.�|��|�w؍Ilu�s�䭏x�#o���:�]�_��'l,�
�M#cɺ�+mv��+2&FA�0���v�jh�@�14�]������U��"�ⅆ�0�q�<�oS����|��cg��B����	D���w�/�aW��������
�#��-�aZ��45����O88y?��8wnj@�q�؛�" �{V�{^�N���n�~�`�<���^N]kkk��N!���x����}��R��<<t�g�����jqlJJr���о�Z�x+2���n���eIq�
D�� E�c�3NM��fWW��;v|l� �Kߦ����u�(�nX˖�o���CJ�R�XY�2�N�o<|����Ttё 3�����@3��� �c�UH��|�MI�#Tc�-�f��#w������1�NV������I����s�Ͷ�U��ᇏ��Yy7(�M̩?��a�*�3�I��O~S-dz˨���J�)WK����
T��}�"�����A��s9jק��4�vIC@�ʁ�SZ\���L׮Q��H��j́����+4��g~˼�\�m�1�Vju50c���93��EP)'o''7>���J�2@Aن�[� JE��~�s�����ݫA�8�o9>:��=]�o�+��l?]��10� ��* P'�ù�Ӑ�W��ȍd���k�8~��P��Ic�����r��G���}[Z�b/��P
�� 9��;9i~^�N�Z�Ĉ��������>Hao����	��ۃ�Ji��Y2	=XW�wþV��q�L|)kS�L~�����9M���pWS�܃:���.��+� ��n��$�8���$�5�`������څ����Jok�
���'8g�w:T�?�Π˝�%j���4���N���F%�:a���ܬ���[^�n8|0O//��(����:(��5N2���3@h�H�;�*����:���a[��s0��Q�GÄ%OφF��g�J����? ����kV��K,��Y � l��	,�o���a816ZqѴ����v���)t�*
ID�hX��j�S�AK݃r���b���n�A���1�+����7@�4����yH�<X{���z���0�g����'rr�P�H������P���vv��߂ ��?_�Fz}��ȻH(3�'�d dñ1m����x��*���Y@�Ђfn�s��ppk�� Q�5�s�����KK�lɴ��׋*U��28S��D��%A��#���~�f�?~���w� ށ������!A��=T�
0�
��8��۞_�/�<7%:��IgC���6�Ɋ�'�x�2^T=ym>��r<::z۴�b���g�e���貇h�j�P����g��KH� ��RU�x��q� ~Z����M�c�
cۜ�+�υp�Gt���6>1V�j}��.}�]=a�I����Uo+���P���qPa :��1+&�~~���PJz��]]ݹ�O3ϑ���箇V��:�����w�! �K>��m^�JVRb1��llo7Yt���6��#�2X;>2���N�|���v�3�Q�[ݴ��Ő��k������H�B=�5eF{cZ�7f~'�b���Vg�^��[��)�/�{��[�'�m7^�[
�JP��<�Df���4j�lt��Ҿ�N�jg��D=�5��>���?��8�bX
X��_����C��b}������ �$k9����l�� W�B��j|_��)~��Q�����Y�ÄG��o�]��-Sa{���&�}X!־��KÕ�vxv�1�3�ԭCo�Q�[Q����Q�L���֏&TM��eٹr#�)0�~�~S����TV��2t��
�h�n�SqB���\TTJ� ���-Jj՜��.����-�C�4�7��D����"K�(����ר7n���X��-�OІm�����@�\\�A�����ly���� M��p��yoooh#U��)�lm(@�
.���t�
���
C�(��2��RΘ��Es�0H:׳��R����03\�]��Ó?>T����: ����3#ğHB�����G����-�k��TkkZ.㣐�AK�W1� ������oCű�'�9;�>&p���:70Ѽ�ϵ��l�u�B7t��I����ڟGx��p�J�:��%x����7��d|�	@�;ЫЎ@�I�K���EfV���I��;a����k�*����. ��������&�(���.w����*� n�pvgk��4G���wS�n��Uᜉ���241Q11�=�
�a,t��p�������&��H�AT�SκIL�]b�c��O2�s.��������H�4�{p��w_�������=?1997��' ��i?�4W���o��Z�%�H��#�?`�jy�<��+P����JaL
��[��*���ӵ��S��Nש���3_�?z��a'��������Rr}����tvwM��mhh�Ʉkk�������yM�1.�L��ӆ.��w�D���R�؍�+�m����%���'P ��6<C�끉}W���з�"��@SS3:]�w͖V�F ����!�XP?��j*��9�΍�c~L>�����m޺�3��ʻ��Z�9�o���_&�-�6+)+O��'���744uudffg8%l@����Q��ķ�6:���WD�\��ep�����6��P�V��R�3T߭��X���y����:Z���a)����5fL���0����8�&�^%̂��
m�9$>��cs?R{�s��V��ON;�����)��@��zQ���)����iv�Pi�2���c���ITT�9��옘�����������c�������l|z?Խ�qYRH���= 2�m�x:1 V�o�PC��$h����u���Z�� E�d�_������񝝽׸��'^�m`�:i��u���h~�t�C�L�?���։?��i�-�~�+�(�~E�JY1��VO���t)��/m׷�&��P`�ꉵ�@��_.�F��r� �.}ئ��o�%�@��@�yk�N:�k��]y�C��������k��0dB|k�6e&��~7sM�����N9 �|9�q�2��ep�ˤl�����w��b?�5.�S�*@\���_�hR3�T�����[L7?������r�pw��D|�����S6?1Qt?pCy���M��|�I��X�f*p3��o���'���1����.p������]��	�'u�ܱ�����3�Y_o��Hl��c9�Ċ��|q�A:��Ί��]���c�{�`rS�P�SMr��ȋ��,ǋ�Ϡ�H�V�!�U �omm������p����:A/���d�y���Q�F6o��`*���ｑ�(�X���dn���������9�}Z�,P`Q��
�� �;��7F�������B<ζ��SRRn�(�������c��%;���ڀ��Vș��Y���6�p��oRp�>Z�@D/���a�kV�frV�;w8ZעWƠ���<f��y��cb�=6��W}Q�M?,8�h�HB�$u:6��3��_x�*���ԤT�6��9��A0���]*�`�T��h�����@�3�r�@�ж(\�f�̪]�!N�bv?�I4���5_���=����v�T�.-��s��1����9?T:
�Wl���5D��k�^Cc#�U���Ufqfff=��fM?�Rg���#�~��lvՎ��՟���t+/��:��G|�o�[���!b'k9}�=�eU=c��j��Jq�c�X������OLOg
552�1�����=$*���K�$���Q�K���)޴�՘/I��sT/:UNUxz$�?�377E�B7��VsTVX��l�jG�������g���sq����[[Em3�sB����:&��7���Q�9�C�@C�p�j9:>V�C����}��h�X`Qf��c����<��Q������ă���\'�4&���������x���ٽ�1��h6�w�ޔ��g~�����߳VU���7w
E\�5اlnn�O��h���@Y�C�Tyi�F<��}�ZY999�l�G���O"��%�+�F�摥cG���T��J~��YBozf<��Ϙ�y���3�qkL��烦��خ������2l��oSxW�f��������LYV����V�%C{���s��s-E{���A+햷�8��s���S�U��3��������+����%�
�''g�R���үb�%���:�f���W#��[NMƃi��z^�8�M�CM����S}��FyAΞ�9�@�|ms`9�ҿ�-8V�^t���Zƽ��Z�K�΀�9Ѐ]9�I���'}+�g֙ŀ���+�f��|_q���*ooG�Z	�..."��\�d��%�3�{�z\-���yҜIݰ��6��$��g�G]���iT� >�n��5����� �yG�I�߿�<�Q��q��z~

=����i�j����7����Zo 9��L��n�_�o?�ӥ
e�Q�?�z0I�G�/��������eGkk+�i�Q�ؒ�їC�[�}K{�4 ,��/�ЦU.H��^gr�{���c�����=�M�T9M�3�ͤf���t����M�7\��j�}5�����a�䰵�uYU�V��
=M�T^~b*�b�6z���/W�gA�y�;��`�'��4z���i��Fa�D����z����˹
��1C������,-����Jf�(��"- )7Vc�����[;�g�g����:�lub!ߣV$ظ�0�z�{��-��&�9'���ΒQ24J�yZt�>��12���;cE���2F�V� @n��Y=	�|($TVS�yu��ЕE�[��ϙ򦁥�:(S[[[�_H�ek[��@��\(&���[��@�Kl凜]wou��!��i�<��w��\vB6B�xn@'��HB����^������b���aV�Uz{�C(�\9���KU��
��+���u��j�|0+�.q/���B�k9�����:݉�!��ϼ��Fr���@���wa���u�a�m~vw���
:ϵc���F<{_P CAA��� �z�8�)h`J�uZ����p2@���u�+ukM[��<�6V���UX��=�J�?�<�)�M�ϟ��@�&����r|���Q�K>�-�i\�B.�"����$�=�	�^~��Dl���,^,�Ie���}��f�|�V\�	�c0��گi���ܦϋ��KoԸ�;�~�Gi^��~�|��Xс;�8 ���Q��� I�Ф9�^>֘���>h��P��ܝ�����F��U�p4��cL���Qٯ_�b�KU�7(����By�:�T2�s�p蛜�w�?����Er=�)3@oAiv�w��D�c@�{n����������x0j�eH�4@��ԋ�ܜYx��묟�ƫ�R�F=c��;D���r	��t6���j-;�q����oҢ����4ϣ�a��U�۹�cS�`Ri�ݗ���� �)|�R��~-W�n�5����(��峺�v���s�%k�"#cc��k\B�l��s.�l�c�8Y��u*�P��.~69�[�U�~S����9�V�d)iiPf ��;*��l�A�//%��-�	��ß���T6�A5K%v���6P����A���ZU焻R.���`�w��^��1��!%�c:9��C�	���CE�T\��rA��ކ�5%�Q2�������vߣ8�?X�`t��*��~���dT|��s���
�CpnJ�bod����z�D���4��$BMB�
�O��S�UM��ߺ��Dn��p�z���籢~pj���K^�NqT��z�	)ݲ�����.z�Ey�辜4˕�k�x�5a����5zU1�$�=<t������XR�L ����̲6ϊ����蟼?G&�WK@IFūA���b�&��F��*��\�m~��~��xQ��-w�o ����ٿ��V���v}Lļ~�w��v;kț����o�:Ď��e�5��@B�7"Q/�h�J3�["�Y��M.��_L�ݮ*u��@6{hp��Td��_�D�Ȕ�ۇ=�������⟘ӟ�*�\"l���J4��a>�ք��mU��G[HaM�j	*�ѽ��_�����34�̪�ǰY��Vm]gb�tk�6� 5��?�_�]�'��^���d-����T���L1wO��Re�.�T�p�K��Wm�;���~��GNp�f2I�����v�t����ᗁ�v���~u������ÒH�ƃ'DE�ָ�%�P]�j��0L�1��~��D7�J�4�y}^rU�wf�}跲�c������˷���z1��\Ͱ=��	�A���BϫV�]F���e�}��m2���-���kcb�V�%���0��3�(�m�4������i��#yM�Pz�������԰0����kվ�*=�j�P���sv98�#�<��O)mW�w]v�G��5��=�\�7�%����<;ޙ�@�4x���C�c��� ڵJ�{KC3����38�B5�rļ9�v�Mf���I�f@Z��k����*��8*��d������1��r*5��0tJ"pbzU�8##��㳛�ț}|��e�w>���@y�?]��/J��Vx~������[[�|�〭A�^��`-/�l�}?�>�@����4��J�߉a�7�#W�ԃ� d�*�V���P�by�~ˈ��~��[%����ܐ�7�z�aA;݌�Ig�W��j��6�ʰ�Ȍf���Ub�gvB)��,]��-h{{n^�!m�ʔ���6����������+��&�K��m��J���K���3��_� �֐���qj�l��9�߈�J��S�����Br��V\����@����i�o	R�����1�{h@�C���������V���gn�E��ۋ�r��_�SǾҸ8���,\�A�}a�W�ȴ����u$йPa49��;�w�)P[�j�4V�;��=�vC�83�d�X$�t��4�m� ���''�

*���JUq�����7�;�����E���n(��n+&I�#0۩~�����>G?�VH�qO����>�
1�?�ׁ�K�R�iv<|"��4�ka"�8��z1&6Q�(EI� K\h(�
�O�GԒ�V�t���K�wrw��z�TIݶ7�ᨋJ��O��Nl�yLOm���w@�x|b��r p�&Wb��4A��0���q�ʕ6�2X�����t���@jL@Hkjj����V3����ѱ�O&�.�(�Ǯ"f��t%"�ľӊZ	�?'�b=�3����+�3G!ۼ�ڭ�Ɏ�S�c���1m�Pxm��cgg�5Lw}%~
���}f��Ѧ�;����iU[�Y���v����?A`p����C��;8L��U0��ƮC�rzz魭-xU�_��}9�o� ����2u �B���h�k�x�����`�D�//�5G�{���bR�XG�)��i��p�f� ��F�����*w2_��ZUg�8�Z��� owv�~]s�����G�EZP
�����&D_	���϶^��R�;���?A��7�|_��Q��<����Q���W�cp˻}��w�Ӛ���@R\#������ ��C��(��zc�||v�z��C��R���7�T��z�1_C��^����7wϯe��3N���[��w5Zι��Ҋ�A6���(��<����{�H
�&�7��:��O�/XR��� ���ŋ��A��&Y��?�҂<�7ea�>jr�i.�� T.b���O��q���y���4#$$,���pa� ������<)��ќ�o�m˞�6d�ui����R�xM�~�@+���%��"���t�>�V�/�lŗ���Lڶ���n���]�R�y�g;kj;n:�E�c�Ꮵ;O�Sé*��ٕ�|��k��t2n�sH��Y�W�tݔCf����.ccTž8�#%
���u����x�k�μ���Ey�O�_w��կ�Pl��;J"x���[(��6ǳ���?�r7���'g����ߘ��m�93���L�-;�؆�ӧOߨ�zušZ���)_��bzܝ�r("	c�-�#�W���sg{��^9�Zv��-RRRBF5��XkC#�����j9�����F�P*1[*���bS_��0�ޠ@�m����L��fr ljjj��g��uj��&�������c��lpn������_Q܃g��Ni�d�T���j}֓sC� ������k��S=O{��"O��P�msZ-�H;��n�1o�)o�I�53^ll,C�
#9>���e&�RY�gƲ��{7%ɲ�PK:��t�J)���uT+�h�OM���AC��U�~��m�������kW��֖_@ ��/��#�O�/E�\E���:&H(��\��>I,��UQ���Y��Ls(�=��J�R�������i�\�M�Y�~��e���A��~�t�6�!%�L鎂��vz��g�m�u��mCرv��T�`��2m��`�5۾�+��1P0�1��� ~O�f�C�+�*�H����V�n5+"�a�e��F�+z��]�ӹ0�X�Q˾�@`wA��n�Tc�͉�!��-�ҕz� aI�\O�������Q��ks�\$�T����b�<=��ʺ���~r�/Mŝ�bV̉��n�ڢ�ĳ��Ӷ�y�ć���?-�Ҿ���W�.p'|�{�;xCt"�$L��r�<ԋ�~��\��N�~��hy]�g��A}���o�����a�s�3�n%2b4x���7Zg�665�ttZ���O�#}���(���/��R�f�!h�~t[^g=B��d�'��_ؾ�L*�}>Y����0~�┑9���X�YE*�KO���-�_��UFK���������pS�"����204�98��Y1i��q�vh��Ko2%�<��=�An=�� 1�˖�i��f���0l"C��]F��:�g���9�К�>{�7�$~�	cA!i�e�<iT�i0�p�!�I�pO�Q��x%�'�2k���զ��$�R�YxVz�����
BV2O^��PS��Y4Mp�T��7�q�{�,�od��fTIiT9�$�-م�A�v�mUeˋ,��^��`ꏞ�����.{�`NF%������y���z��o�1]��#��"����9IhB�»S�S
�I>�%�u��A+���9��f���2O^��˻ h0��V�nX<�D���o�
�Ka^�ċ1����>I�{WX)�ݬ=�]���^z��O�w��}���q��!o�fƵ���b�"�τ!��ymy�-���� >�*�W�X9r��e�����\E�i�\-)�_|����>������=�5����ig2�z/���:�1��+O~la57E{�JT�]�sX�/ ������:�>W�vW����Mے��
�`V�<'.��������Kw�����m��&��xF��2��J�zJ���]N���N-@��0�����|?���#ؗ.ELp��;O5e5�[�Z.���".:�I�
��:<=�{G��:��p7#��`>[צ�X�_h<��˲k;��RG�x&.pA�]�U䎽�Ӫ�������c_'����M뼊dV�s(ܼ���(��f�a�>�Jmd�Ã�!}��m&�t�	�ӷO���e��'�uu'���,��������f�b�_T]'�A���@��l���I]N��x�y�'���
gN�u�����wI[^^�o杻���ΐ��v�>��j�VY㘭���=��c�Yu��nAU��C��.Ů-��[�n���K3��Z���0d���E���M�>�/��T�ݐ+�#���DKg=)��ʱ���00���ĥ!��km��8�m��=�B���^h��=�}������)�ﺦ��e>��M�T�4��x�H�_X���#�=1|����?yZ���H˂9ʲ��.*b���z�H[[[��
��0A����0Ѹ���>�ّFˢM�u�n�F6�����w
��,F� q�ɻӁ�C~���13c�,b[!{�|
���~�]���Җ������)ACG�zZ������o���b�Aھ�uӲ��҅��=QQ�M\���G2_�hlo#7|%v�]Ò'�{f���Zt�I��L�����p/DW�V��E٠���ǟi,[`�;��<�i�#ɚÝtg�����i��b�O'��6C�����Vr�ӣj�-�H����R��Y[c� ��:������J���������Ғ܏�_S�Y/ϖn����V�)fWZkpg�������ݶŶ���  ����<q	}_s����
�tɨV���)J�'��|�{�9Ue�(	.���8G�d �)f�?��� هl�v����{r�`�Y쮖K�x!��H���Q<p����%���ka��)������;-��C��M�^t�|�� ��G3��aJ�&��b��H��j����p���3nv�7���$��г}�l�5or(��6��_`X"�B=ww�ellL}�v��23���Y����c��O+�i�@z^�}�ЫĿE����-ڀ?=8/i��nɼ5�tww�g�.�$t���cCKC�� P�"�R�9�Q�G[��I�^�z�Sqzyq�H�ENqߔ��(�Θ�Z�V*����(�\�ş$U��-!k�����ڑ�d����7�.*����X)��+�4̜�j/Q�
� ��ҏ�Ҳ$?�ׇ�0;5��M�ԛ�`��'���V�R�-љGeT�+[p{BlU}Rчe��m��n|�H^��J��O}S^�(��O�\vZ�����I��r#�֣p��i�6��ٿ�C��?qJ7)�{X���y��}�����*�=˕��n�w��H�84ivA��x_�d�=�rH�g�4���j�!4iqþ|�/$$t4��Ԧw�I�݂w�6��D=N�Wf�?9q�����x�/��5��2~ϓ"VE��󇎎j&Z���������j
�6ۻ���.q.LFd�2a��Z|���_��
p,�Q�Rt{�Z��w���{r<cn̸~&gܼ�[�Ўݏ���S۶w��%?z�	J��[_�q�_��d�h[c\T�y�q�`a�T���)
��!�x81e����B�|>��an��#�-�#�z���pU�ez=Fا_�m�ުZCwAw���r|�Iد yȑ6[I|��c�>ߎ��}G���n�3j��zOOE�J�Y���J�U=/�4���A��|�b����>%=n�������RVVnv[��2����d�.Ցʒk1Y�R���3�#��(�^z	1x���,a�J��x7v@v���$�.�2��}��M ؅��
EZ@sI�O�1nZ{o'�ƿZu�n�E��@B/��mX4�E���X���c���ؤ�� yY΀#i�,'����4��|�$�Ik��1b2BsW�HR�
4�5��Y��a����٦�5�"	�}/�H>fA?�H^�\��l;tz���?�6�u8�������p�gMz̚ԣ|�#��v�-���{b������������~p4��yUj�{�^��x��;9;���9�
�H3����ē������Y ���O��>y��	:R�����tz��YͰR5��K__�
k�ͨ��E���~�V�]�	ь_p���,�LT�@�t�m�B�*n�I��0���-Mw�88��q���Q�V���Q�^7���<��Jw��v�������P�?}ɋ�in�e� Ģ�"�05�U+�۟�����=�� �FC[h�MMM�P_�%��=�H�t�P����`t=6km#y9�@��o
צf��T4�KWQ]��ӐU-� ����b%j��B¹��[�Ehq�bTX1���� t���sIO�kҝ�.��� Q�OJ*|�	/N��v��M#���bE@P��j���i�Ċ��{�z��M-6J���Ñ�8���F+3���i9�ݺBL���������M%�o��%`��wc�}6:n�����e�Fm�`G��0�e��ý=�_�>%����Ҟy�R�~����$�Y���ݾ�5hn��m?���q<ck?[����������9
0�e���cwZ�p������X��1/]�>�$CL�8���w�4��K���3�ݕ����S���2�����#Tsgc;F�N�-MP*=�R���S�hr�ѫ?B���ho�5h���Y�1ߵ�ӥE�'Ѝ�h}�[?e���#�@K<�H��S�.����g��~�w�l�4H�[	Dd����ѝ�x�qy�JF	������4���w�f��o"��4��J��v-�5w|��mN� �� ������{Z8z�̽�a�������E����R� }��=�qooO���N܍��»��l��K	RDh r���Ax����-.jݩu��_�Z�fIF��w\�u�+9ő�4�wo��D�����T��]K����F�+־���4r$���T����L�f�z��~�bbܦ�] ����p���qC�ZbACMU3�(��Qc������F�%�i�i��~�◔�`���ˋ�0ͳ����Y������;��A{��kǙ�;˧��`����E)�jA�J���,wq�j�k��t7p�3��)RA���V���'E���6	�g;]	�KPa#�	������*+m��#R͝�F��U.HU�2a���F ��47�G߈ ���;y���Vm�woe�m��4ޏFS0"���~�ES�<¶jSS�k��Ѯ«��)������9(2���$��`i��}'_q���M����"wp���ʟ���hoTX�����|��J_������l[���~������ ��M�Շ��P�|���B�C?:�ٟ��V��/9eq>.�-���ͤ@F�+��wz�:�P�����9�y.�L�S�]>��0u/:�o���R��� �p&̞��.�r͕�a��l���u�)<ok�G�Q|��]ϙTzQ8�w�=_D�A����.c�呋�P����a��t��y�Yr�L�q��L���/_nX>����3���L�0ē��4��*K/��:55F�� ����m�Y3�.��&�;&D�|��������s��',ͱ�5!���j������������^]~c?�/j=Ԫ����^o0uR�Ļq��5?��J3�p���\���~Xo�l���M�R��Dl�GX��#��q�܉�g)��pzG

5
�jy�v��a�3
�5r$���i���vO���H��b�JF�e�>�����X��~��ٶ�}K��4��c�9���CԔ����wQ�)@#66� �<�MJJҘh�Im6G8>��Z�Am|{�*1��6+9ײ���F�^��ZMK�u 
����=�S����~�;	]�G���﯑��Aሔ.��*vr� ���@���<a��0�(����~>?w�k��'%�?*Xͪ>}��gAp��޷��#8n�h��z�$�/�5��������S��۲�L�#dI���.e�p{^Ua)���y��#��4;x���㛃>�]�m�?��@���*����O�11�7A��k٨�&���YZZ���ׯ�@����;���5w���5��VcdO���Nf=o�4������p��7�/��7�m��Ode��UF�(a�h�=�2a�~�<p[���r�|�*�������.�]O�t��Ԯ#�q��rȤ�0��0�Q��/O�ʋL䬣XP�/`|�J�g1�����90�7G;!P N�����#%N7�-�{P&_c�\��p�|β��1�e�Bg_K�k@*@S��k5k�bJT����"+�����-xp�rW0K�q�� �'E���Z����ڑ��S��࿋�3����A
0/�gN6
�s�~�ʇ� �T�+e��yX�=:���&���C{+9)a�&ME��A�p� ��@,�����#a�	~����^"�����0�b]��$5�t�I�q^�����ˑ_�4,�@��q&�{L�����1{yNp�"-���R,�4��^e�ؕ��("�u8pv��0E����ɗ@v�n���y��f?�$W��7x��-��(n6�z�ߴ�ϭ�܄!�[����l�C�ڒ��[^�Y��G<9�:g 3jk�cT��d%��X3�m��M]Pߺ/���d�����9b^���[QU���w��4��	��r�X|B؛�L�]*4A��.�)��W��=U+o#nǸ�?z�)��4�������S�p�ga�z� �ג�%�:Q~o �j���s �,�f�"D�4����p��S�a��dI�l���N���6�~4v��+i���l�ͱ�d;:��jB��0�P��h�6�D�ڌ�ӱ��z7Ě`#�y�j:;��c;���9EU/	-	K��k��91��9u� Q�0�q7@�	E��?&`�ilaD�%��2����[��H�)g�铙��Kǽ[��t)C�ϗ��S�c�d�����ƞ\aw��*����K�s�.����]�a�����	�	����9�u1=-��O �H��2v�_���F#S�	c�[��%T."#�2�v�{:߿��syq�;���9	�[EU���eo���,�����\X�I4��x_�K�Ձ���	�my�Y5B��XY��x�qw6?8�C8�=uF �����j���|_C���_a��D�S�Σ���E�7�r�|��rn�㜻�?a�g�)��E�]��2NAUw[����������3�WӦ���W�檛}�G�mr��7���p��2��mghy5E[	� 5%�!"��}��]�bͫ�.<�}S�5�����-���M:ڿ!�q14�&��
�"�S'UG�.��zwl�n��a�<$d!?#����Y����`z�5����E�����O�j������)���=|S�O{��v��Q������0��u\`�a���/1ȓ�F�y��J����O�rް:E���&�{*�bee���A��窷�B=����6��� ��-����0˥n�-�������Ĩ��KMF?8�C!��S�^�~�Ǒ	L�����둙5�l�l��(��[�M?3Og���[�l��~�wr/F?���D��\M�\,�i�<yZ�=�- �m]�{���p5L嗐:ޔ�ì��88ǘ�ࢧ�*1�%2$��夁S���kl%K:rjqZ�#=�[3`��_VD���ԡ7A|u�����#��Qү�o�]!?YO=��LH���R�7\�3���s��,I��ȕ	N����u���Fo'^��:'����miȎY�?�A�Hݜ
E:���/����q8y��K��.�iW�8C��5�������Wܼ������W��_�x�vǹ���.��ȟ
ʊ�7�F�/s�����\�A�_��V�/�8)c�c�%<��}��@s�S�_����?�aA�T��w��j�X�����9o��>���h3�r|O�Ry󟼳݅��j��x��KF�*�1���n�I,ݿC"�w�jM��KL��1k裠j�%A��| Ճpo���dbbz?a��{��d
'Mu�:�v=-����y�Up���Be���_ǡ��Q�X;gPԐq��9}�t���N1��qȣg@��#�� �E������Zn��=4L�G�z��9z�R;U/"��"=���	��(wFg� ��X�mX|_�6�{��B} #��y���������G�0�cX��p/���Oռ�iܩP�oݥT$����� X�!+�+����qj�4����������1���8�jÚ0�,_"�R���K������^�b�Y'u�6g���d�
+������p��}�Ju�� 'g��+}q����57w�9��(��)!�}/gE��,@�Wa�M��9�(�h����
����mA��PB��.IA:EJ��;	�Nii�.�����f����{ν߿��yD�k���;��c���n�P�V���j|�f�Q�3o��[��n�5Q��)���R��fM.|��=`H��nŘ�t"���4 ��*�|�G��Ls,�>�݋[�7��GQ���*��*�tO�Տ
����|D���K��9/��/�?�`;Ra�'.�P�ޗ�D���iJ�p}������c�_J���-��rw-���sn�T*��z|�[��}9cj����OP�ж繋�Uo�:�8�A��y�İP_)�,"	I]3��4d+�����nA�D�G��X�`tr�����_f��~ڔIs����BY(u�t,�%��Z��m*-�-)�Z~|~ך�H9������U��9�,E>��r8K)>�l��H��Gt�=�L(?!&)�����+P9Ej��,�����tZwF���^��B����A|��P�r��G�����Nd�n}��B�l%֒c߬�;鈙jqFҎ_FOA�E~��cR��x*�~�2b�nt��@�	�N��ӻ���k���X�
zlu�goh�V�A��I����{|e������Ajʾ�D�A�~D3���+M�E�3S����AO���m%�Zƹ����y�U$���ʋ���/7^�"��5 \�!:�*v�C� # �����;�*{V�;��%z�<�i����{�F��0&����E��'KQ"�����r'��1�'^����T���!"�6F����bxg��h�ɿ<Q�9��:�����J��%��X���̋�̋
ĩx���m|i\�G9�+9����ɪ�b�5߬�����OD@_��YJ�1�7��!�W?L�Nի:k	�g"�S�Ey,X7�֝�-�Z�g��;��1)+18��QP�q�^�+��j�\���w��P�O��5�����^��!m;�/,,��N�Y.#]:+'�<�g���I��7eQ�o���������,�0���R��l��`���Y*�F��e���󓮷��Ϲ�;o����p	m�u΍�8�#h�v&8)�����rB��Q��dkR��Sw�D�b������|�jM�Oj:!+�{F�����]��uv�f�_���ʨ��$�`S{d������#�v��X?LF�2�y^�z]�	(����ῂ�-NN$3�S]=}N%V���x� r�h��sN�4p3?h|��P��0恡����!�H�!��K���$�i
�ܝ��]����	�WfL��L�2]�9��=%�R�Z0>)#�R�S��䈼�{П��Bo]%u�Ͱ����8���wS�
��r���(���e$���p'�4oBV�/�X�6̼����{�>���`����6�3��M.���y_Jo�?-TB�1`F}����w�=~�|\q�9�&��B�B�HK�y����w��,>�Ǐ���irˏ{�}��[I���h�ŗ��~P�ex��"�]�����{|}�z]h��55E�o-Z�o�[����C�nP ʫ���Mȣ?iqpz��z��f���hJ�a*r}ٝ��@o���W����r�6m����9
+��)�$c+Ϡٟ�4�5�Va}Bq"��E$��Ե�&jf`�u�;���6ǌ#�SE��v��������l���]J�ٓ���hs^�]ى�Vz��Jd�N:�#�Z�GR�@�Z7�q�}K���������-U�bQz��$>���yK`\=�|w!��?��[/�(������E��S-��H����q���M�.�[Jl��yq�g�m^�xw��rr�l�B)�Q���鞢�ڬY���7?��H}c�U�.�n7ts�%�{з�[���J����b������i~��=�?�ٍ���'�"h�9�����m_�?o�񛴚�tR5�ҼY�i'Y�T��[-a�G�}�{�CN4�y�	��^���0���CAz�l�з[�q�����M�j�0�\䲋�-r1�܁3I�᧔�f�ժg����Ab����x�OH!8~��|�B���Rj]&\>w8ؠ�g��t��L��ֲ�6-����ѦxiQ��o��˺oM��Y#Qb7H�f��y����Ӕ~�k`���&��F�^6���:����#�C� ��- �\T��u��66e�Jq_���|�cT~g_0��}>L�e�*sX�m-4.k%�!����V�f7�l}���	f�ͨqy�����������R�g-�L���d_���˖���|R ��zw#� �y��Qv��]/߅�q�M*'�S����W�d���F�*��_�А.�ݘ��}aƻ6n;}H�����1∯A:@Aam�<́�&�{;tXd�%��s�����{�ƹa���9��X�4�cr�+��e�~�@Zc��ZL�鼝P����}q��;%*5��\:��'�4��*����J�����mٹ�� �t�i=t�_B��*����L����$�����O]q���! !�*$��{�qu�H��&B�sU���|�����V�1���*�l�I܏���_�����zC���S9x��I�����3`�Jy ��V�~ŜL\x���껵�sQF�>���
�P� ��["��i�H@�:@��� ���ok�M�[cߺ	F^(����5��Y�?��D�mlI_�joOw|dܭ��yY��A�[9�nC~�=��R�,��b�rcIf��##8999o4���n�^��o��~��-r3��B�|r;LZ�ݾ�8x[� #��1�#Q���t�*e�_�7��D��Vm9ݽY�'�C�g��+�wǟ�`W��0�o�NTy��s�7jp��`ﭷ��ك�򞅄�9]���b���f�����"[��y�f��ܭ�&{<�J�� ��Z�>�+3�,<!	���ߐL�<=͗?��� b����kk�%�ߩY�(�[���6(��^z��Ͽ<#�G����|�Ԝc�?�������Q���f�?{�6L���ð��
�G�D>��+�Lh�n��ў����֜�s���<�����������0�%>g��V��g�FFjot�`޿�����bB#ꓺ��1y��v1���)?�7x�yx�L�:���������#MM͟�~��L��"�jHd��]P���32Ύbb��>��Dj��֜A$�[j���>|��ya���]�
WW�.���O�s�|��i���QZ���L%�_���\'�*1�7*F�vu�͊:��o���`X�+]#>)�ml���s��X�ak�
��Uצ��T��_g��Fc8-_R����8ߘ3<Os���0�K��_�
6��4���]~+]�hh	oO=���9��G�}�A�n��d5$fܲ�����s��e~���I��-�a�^L��ubb�>�@�/����.$��پ1z����^�����0�!���'��\�x�n�h��x�u��O�ש~m�Zu��gл����&bA/�%�n���ޛn�u������x�� �K#�{W��~��9�� ��)j^��P��^fz�Q� �t`����b�d�$��]�����Ꝁ(��[cI=�>�>�`È���-�\�5�j�u�&�h�߫�y�.�R�������1��0�O~�?�vUa�ɢ�}�l����П|��5$�Y���ǩ���Z����a���l7�Wmyll�1��u���Ʉl&8
/J�B
��K�Z�N
���ОM1�C��8=�N���*�*e@1'66����L~����'����v�d��J��<�9�)�OR�F.�/$��&�2>CF��ZU��;���W�]GE1,��ג�����Vc@qJՍ�i�H��|*�����;ґ�F-6��27���$	�Z_<���r8o�=���L|����)|�O��F���f�ל9��Ny6[^^�ފ%�5)?�իW- ]c��ic�]u�^}�j��9�+�|�	~�E�_A��o�,)�M������'$�N�|9e���C
'�Ϙ:6�V���ԏ3�~Nj�z�Pj>2�'�����5�ϳk��WR�}3��++��J oD�;J���A�+�$�S����
ȗ�ΆJ��û��̓�>Zك[Q�)F�o�ghk{�fl�_�␑��A1��?��)�sl�� nˇD%��Rk��ʒ�͚=���%;�O�.7�D�\Z���A��Cg��q�Z�����̎;��^�_v���~5��n?�����tHuq�s-����2��bTxVkͯ�fه���5���4���ȷ��GR�(�+;�ʕ��(D��1J=��ǲ�g�U�9�.Pl���?$*/�ǆN�~Wk��fY�>��.:����^��F�_Ϭ��Y]�85� W���η�8 \I�,'�Ő#_��j��r��C��-�}����a�=����/F~��Sf�$�~/�y�����; %R��D�qӝ�k�����U��PO�Lb��p�{�wB�J��. v�φ����て�=흃�w���������J?g�н����Sa�a������ѿ,&#V�����0���f, '~}�`�8�)/�8 jV��.>���vz@:���[�{���㷭~�[ʑ
C��'@�P	�?�K?�~Hw}V��k�h�c��zy��u+����c��ϻ��U
TUhq����,��F��oo����$;|�����l����/ip�E��qh�Iݴ|�լP�����z��r����C>
"6iQ���g�q�>G{�w}��u���E����	ԣ1$4t��.ue�;P�!lU�� �F�t�<�u^�FݟU�ޕ~��\��YJϲ�M�_��;} �:d!�k�X�O���:�(
ɓ��A�<(Yf��x�/��Y���ͽ��_���P�����u쫻~\���	��͗GVל�����m-���n���A��������jam9��L�a瘐'���H���5+�{����8&ݎ��@��ϝ��K&��r����[��E��OŰ;�=\��X3���?v�M.��������0�~�հ+4y��Ed�f�'Q]o,-�߾s4 @���
�Yz�1a�� زR�-�XVV���;`�3o )�&�/�Է��㣥:�=ҧ�/O|�O�ؾ��Ea���b>������E��_��ϋ$<A�c���he�F�w�nB��98
�� cvW�%�'�������TH]�|[�\�g�.
:�r�����Df�+��8�<���Ӌ{mn�T�E�{�h��� ������<��x��)诖�ުW�M�� }(��q�?3Z��}|BpWp`����Se��fBwۘ�VU�K		��?��<	��SA�v0�N}���nZ��h���C/����[:�� &o�|�*y�o|���������v��k��_�&���P�w�P�}O�A��@?�,=��V�L��o��m���
-��ܽ��ݰ������`�N�ZX|��s!g{���Н����9%���_�KK�iAؕt%����n���tJ��9I�9%�h%����j� ,�+���f>��ф�����@��L� d��.+$��<3�4A>/�ߺ��m;���QY�FT�ڶn?�Ǘ�$����DD�?s�������KS��/�۽����Ĝ9��Ey���%���>C <,,,��#��O���8��'�ֿ�8��"���� �HuF���>�Ըu�Faq�c�r}�L�n��A�kk9�F�y+����T�ҩ��gAF�m�`C�$��Z�}�{�e{y� �X�`?�DUiSShQ�\����4ϳg�4xxx�/(��� ��o�߷��T���r�IZ7n�6Z�-E��Q_#�[m����]����t�M_όg2d�GV5�s���ǌ��4�+Փ�v_J������������洈�����:�N��d�� ���	߼���,!��ܶ���B��h9�Pp��ÿ�{�N�5�j�-�?m��\ku ��Ѩѳ�S��v6���fG��l?��M�ɻ��ܚ�U������ 
�dg��1���U�������-7���U�Tj�M�u�[���brb2�'l}��4���X�z0�����8�U�i*
�~n5e�L��NQQ
7��z��@�؂ss��7
뛛�e֩��J�'-�)��󥷶����o	�>ʮ
TN�9ٕ�v`�sKQI��n�<k���՗���oa�3��	yƅ��Yx��Pi�t����S�j�;m�#�Ù�����.�_���hj$�ߓ�����}��2>!Q4+���s)�#-����P}��OB����߀m���F�to�ȕ��)i<J�㩬�;���C�������/��mm����]����������qX��dd%K����?�����PTW'w�D��4?�V`��CS3��Ǆ����~U�|/<�c��������O�C����WQS3�np��G�k�4��"Џ�m�"3��~��
oߔl%���9(���f
N�:X�'�:ɼ�m�)#^�4y���G�%`�:9�AEE]��^�O�%l��IIIQ��4{ Z�{=��?<x'[DE���ӿ��$#*ټ�֯N����0P�]���c�����[Ӎ�/� {�ʃ��\t�grnd�r�p�y�U]�o�-0g��2F��R�ƠWg�ƿ�"<�~�ܜ�Jf2a�	U(�
ϡ�)�����PM�u�]xś2���DEQ�I��|��pܤ,���F]�x�]S��t`i�OI�x�����)�ŭi�&czP�����"y,wE����q2�є���#yʶ�Z��5��tt��ө��V9Q�׸O9��jsE��%�ћ����>o~?Ӆ�6������7_�iV�+��޾�N�R���.7p��Y9��~���� 	���ò�e����'�t��̀n�B@�~j!�4�V���@ �?%��Tڰ��%TǪ��c��PV��roB"��%�~�k�vQ�3���&�(���r�9�f�Ak��/G�N$��y={��|�w�;"�38������d�C�{ֲt��d�"�^2u-��55�D��n��L�K�s�ԁ[�����(=���[���hQ��F��ߤ� !qty�sN�+ǯ���|�<�R��ow��m-ҾB�A>�^�,۶�P�Ϯ��p�l���)tT����~���P�Mm���D!/O;v..��4�XFĚ�ģ��=����8Y8>UD���}��k.�+h^���e�9�Ɉ��]+�<i��:�%P�X3��F�"g�P������r*��6�2GX����fҤ%p<�����U�Mî����{���Q�ǋ�C�_I^���*�����!�V�i��h���kn����ds�d����,X�h���_���I��z�óU�`�\��X�9�mS� �����T;*�A����*2ى7J���ZT����@ l����/ϏW���ע%�N�`]�E��hh��Pě�������-Gd���^?�j��~v
>�6yN���Z�KRN�i7h�T����]tvvF/)Stx�W^�u�v��4���o���
u���F؟e;��{����B� WLMMm9w�.���J�̛�U44X,�?uHj�����o� �W�V��`vS�oh��Xt*Z����^�xdU���a�1;��ym�+Jy��T$ZK)��P�9`��[p�J=M�$�Ϻ�}>Ł����Y{����3=%��Ca�@y�������Z��,���MoOՏNM�T�j3�-��$!~�ў�j��hOF�d�c�<Y:��8h��p��6���m�&��B4��G�{��6t5��1:&��5���gN��w�c���k	d~u@��p��Ҷ~
Ec�]���.�99QQQ����f��!�U�/_f��d2�"[o�x p%����@��F�s*�L�#�'����4!�p�C�yu��m��e��$��n����wX�I��ן��vAi��,MEZ�C>b�Ps$38�(޳s���1̎����
��:�I��x>�b�Jy#�yϵG�h���b�P.H�u.���p�����T�[�⺍�j��Gͩ�KG���N��^��Ed�	���k�����Fv�%�Y���Ծ9 �LMT��o�6@ܤ�ك.��W,��0+v���Q~N���1��/�&F{]�o����p��&����G��s�	�'���:6�ݎ�<���ۡ��#�
PJ��$4:���A�p���z~Pf�)��c���f#��&��/��>)�`�=�|���)��r����u{��PY�j6V���1N�Bg����|��]���ڭ
�������I�z��ı�8�ס����D���ͼ˞�z��������^FO�I��pbB
Vt=��&���H�_ϋ���􈃟���̵`A�HSSS.	k����<���9I���==�	C�R�{���DYR�~��3����-���xH���Ϗ��@Hٝ��V��(-�N�O1�<�$.��&�sMM>3K���z��X����.f�+�b��N��<6�o�ҝ�Bw^@7�A�i�e�U�L�������{���+tbד�����S��4uX��C�A�\n�AUTW2̢||dr2�Œ���FL�N����w�J�c�<�",�����Q��o	��C~f��g�xA+�Z�3I�lb�Ka̰:5�1���8qC%X��絍���cR�ۄd�?)v�n,��,^��,i9���o"Oe4K�Y�a�QTEE0��6 ""RQV#�����Dz�g��$�|UUUt?�Opʀʟ�ϾQ��%�P�^z'm�i��^�zt���G��i׿�7_Psf-.~�l}��4��2�G�g{�Kc���h���/�k+� ~;FE��S��ϡ鵍�њ])�nk�Z�3�?�a/��� ?��r��A�+ �!�556��+'g��T��-~���s:)++�����%�;���1�]�#�u�zrkd���Z���_&����Y"zAɓ��0q�m��E�v���P9z���t����z~�3��Sn�v�E��`��t?�R�S�9�\�PK&�%%��I������$���=��嘘<J�Q(�z�$�<k��rHN�h����
�������*��i�-�%�c7�^^ƀ�ë��� U���hm/peI=��
''�Tn���9y'�,�a&�0�AU=�b�����zw���|���\�t��7�Z���"Ǹ�^d��u>���?���p��9󃠤�ht}���ŭ� 2P�T�B�aP1:�S"@۠n���5/릅rD#^Sa�����J��ċ����tGC����ń%�Zg7!���m������2M�F�"S�z��:5��7��ǽm�NiF#����m&e�F-o-��qu}�Wx���M_vrHH�1�y bҭٞB=�����b��.ڌ�cړt3_+�}N�hEhY�h�$�W*��g��:|��k���^j�8��c���0�/��'p��M��C3�!S�+��J�#�(�zkG1�Q�xB��Hm�E�khIO�c�-�R���լf���m�\����>��s=]��'����`��U;U����ή?�~i���(L7���|1 ;�^/��E�g�p�O��8o꨺�X(Y����*�� P�?�z���E�V�҂��L����>u��։(����%%+#c���!����os��KaG$
;����u�M�����ɒ�@*S��c�˘�i��^��mtW���8�~Kq=*)�$r�$q���F�,�<Qm��O�D����O� ��0Κ{P7e9:2b�~��S�h/�¾a<�4�(��U�fRƙ|OA�cS7r��+Xu��R>��B1�4~h(㏊�yyRrF���0~RX��c�L�(<D����ol��6�½۱��&U����G�����:�	i�P�n`�����W��Z�0w�ɕ�R0������ԋ��vӁI�)Uf$��x����L�d��h�=��	��ѥ��K�����k|B�n���Im���+�H�9ئ1p�o~P�rG����F����B#�\0Kv@��f|(��Uǵ�H:!��{��2���ɪ�|�SA����}�2r��-��i�B�_
e��T<%t.R#�_��%Y�I��u��PZ�%�� ����=��t�?�n�j��s!��J��Ǭa�j0|@����<�=�3ك���r���ɩ��a���<P��q��-+�[;����h����
��t�����j���^"�PR�d���diZ���O^��L�z�^NXޞ�5>>Um��M�b&�U/�gB�v�׈������u�p��X����<�X�4IrW�bb���J����T75	f��x����53�B��h�c+�N{���cC���-��ص�\&_�9²Z3N�1��~��A�N�ӧO./4��9���cc9��v3߅�J�o�N7���re�|�t�u7�um����8��:z��[K�<wI���e���K��rD��fv�Y�03�:�b��SP���'���u�iG��= �G�~A���8Ƿj�CuTU��'���m�N&ܟX��Z9v�с$):3��d�s�6��$I#?�?��]�>���ߨL�Wײ�S+|�n�۵D;3<e	�8=���GDBͫ�nE*�c"w~f���lT���}]��D��4G���+�uf�6��:�������.d�����j[���;������c>���,.fAe$Ń�����6ϔ(�ʥx<�?vs������,	 6 �R�g��B�?�J��m;J�j����ōG��FUm��]dx�8��W������f
�V��P�w��u�b�qGP�7�=<�+T��H��ίG�'FB�b�ފ�ۚ�M��f(!Ǳ�?��쥤��U[�^h(V_�G�G% �?9y~II5o�>�J&W�<[�ccc���ܙIN���nz}��n������/៊���(��,%.�%�P�}�P[{�f�A��_����RRW�մ������4�x����p��~}���Ծ�Nz�[��e���=$or�Z��N&'[�Xh6�L�!��D.sd 
.�&��*�)ccE�����F��~4�e,}�x�\�20�t��B�f�<'���G�>{�5�ړ=h(N8B�ɸ��'᨞��V'�!�[�����R�Jt���/�r2�+�����&�<�)��D��|0]4 gjT�ֶ$�����Y�0_]�3��$��$�?��Т���- ��@}�F�u-�-vF��ʚ�n*݋o6��U�O��p��%Ѫ�Z92�{��'��-�^?�Ǎ0}64Ð��˜���2\�;�?p���"�-�&&&,���J�װ�]p���J���>���A�Z���S1��R��Me�館4������ 5�#ZK�߳�{��� O����t3Z���`����ju�8�����q`�;�.+�Nr9`�����r�0"]��!��y:mҒ���BA}�q(�̿h�D���~�}=��Uo������E�Lj�K0�2�{0'�1
�G6�e�a�b��n%�^W.��=HLNN޿��w���y.��\��-%ؙ���:c2T�4�~���`����u���(-gy��Hz8��r}��(^$��c�d�l|����oky�VW8/�o���~JA��^�\> Y�
֒��v�ڑC{_�5�rٿJެ�e���&�u�V9n�����v�ceu5�c�%e�����ˣ	�y��A/P��Ō�#?��hN��G�;sGm���� !�}S����������saBN��<d�Q���{�o�A`j�~��h���B@@`}s�w<R�(NR��w�����xy�9�M��#hj2W�����{�{���?��) ��~����a?-ud5x�o��3Ivǹ���K��5fe�0��)Ǥ�B��A�	l�Cm]��f��oB����S�Ǹ������g+P9uo����ļmq�=5���޲㌣?J�>�%%�P��d�3`m�&�S��5{�����V��"A�vU*jk?���J"NEB�~12hu`DTY=���F��CRN��eC�&�$Y�S���mm�����=X8��<�0�3W���X�
>_�ݳ�s[,�w
��@0������ث�e��v}(r> ӳݎ�� ����F��2�r����P�����&SC�}y3jy4�h�~f�'>ઈ��ENC~�TF�2�r�]�����ӽt
�C��p2n�Z����@�ä��$���UϷ]#�{6��Z-�p��+��KX6�	�	�p୭H-�_Y�f�:��a�J�d������?磀'���D�����T	#�������8-�J�:m��:N׶���܁����W�U�i�e��E���:M����?���*���!��V�I=���VvSSh+�Ϯ��	0�H�S���{���9���SQ]�e)z�0��5���lg�ˉ���	2��6Mu怭6�E2��4��c�BJ^�~�a��f�Roj�aKޠ��*��/���M������,��x!����9�{~�� ���p\�WݬJ�Z�x�f����É�LQ��kd�3�71�����K�l�N��P�BhGF��X�\ҋ�~'б��2��EB��_r|E�Y�W��#�0�����^Aq]~��5�d�hǧGT)��m��������s&1lx���<�d6ڐi��h�t[��C6 ����	k�|4,c����+	7'��x47j-�y
n���8�"t�%��0���
,���Z�L�X��vz��u(���\���q���g{ˀQ�*=����������^2��5������sv�k�ܶ�]��ܯ����зڷ�;���&����!���ʑ����Gl����ʰ�k�\B�%��y��+�jj�P�R�rM�l{8ƣ��5��~����]��|���v~�n9�k`T�����`�}���*�O%q�(�.�z���ߟ�O�1�e�u?�
�ݩ���� \��b����`3�l^圈؈�%�W�t�_?�d�>�w��������h��s�-�ɼ����	�P���s�ig
�=��ˤ�(��S�'���l�Ar��7r^�l7����ѽEù�	Y�;ѿ��BP��HND?�n�y�ɮa���X,����Ƴ�	b�VvY��ᢹ`\U���o��'�k*'_�ɗ���H4�9y�wY��r���K�u��Db�zX������ݻ�h����&������[��:Y�e�D`_�b��M�K�0����_ǋ��L�
HH�w����"��:osLY��/쏞$#܈HJ��3�<�z(T�5DL��Ie[x�v�&�x2�8���s��J���yyP��z � S-}�I��EI�U�e���{[�:+�׆��V��W���&��,Yw*W�ṠJÓG?�h#�ĕ��A�r�&\�d�dڪ������ o6K��~6���K+�$�P�[��W���<1����X �K�o�w��*���*v�����8�S�(ZJ��Cq8��o��~!}��H����-�Fhn��֣1E��G̓OdP.[��Ժ������������}N����ꂪ*��q�Յ 	%��rF%�`]t��蔡�ў��J �?+EQH�%w�L�q�'�)�9�%M�Q��d]B�8�:�9l�uY�:���o9iV�a�3�T7!>��&G���g�j���(�9`k�?@��%)o_���=�NV��s�o�|K }�,�`C����lc���x@�C�h<׿�˅M"�l�z�2ɹ������)K�u�76~�҈�kT`A[��&��[[}�ǡ��>^O��'(�eߣC�eX1��w�7ӣ?%IRyw�?��%��sQ7�Q$�ht�Ӵ<>����#�����]��p�n>�����"��vގ�n�ԍ?<-�����̫���":D��F�4�����J@T�$�)����"i���%�L���$O/���ᛤ	ֲ���._��n����Q�%ȷ�����]�~��b����_��ղ�e-I��t��,��~�9�W,u.�{�9'�\O��>̷I��?��ke��}u���_j<H�qT�6
��>�C����^'萴K�a��0O�Ϋmń<�9�H
�4�zU�ʶ�J�����H�y41������)/���6���o�N]/��h�8�B��9^}m�a_2x�F��N�
)w�pdQQQ���������
�\Ff2~>n&v�I��a�C�=[u�7�3��Qo/�	��]��?|�-�cX>n�U�1�c wL�TXc^c����X5V [?��	����\�,VɌO4ҫ��h:���3��C��
&�F_6�����O��0(�g���H�ݮo����ڴNz�<֯WbCJsr�}���/�����@���+{��n�.�:(�	�M�~#QQ�9����ϧ�$��V����x�g�E�^[��M�<)r�?(�wZ0{�s`�G�PcyW��	`����.n+2��C���$i�w�r�D��7���3���#6v�<,%�z%bz�ֹz>�ny	�%OM�1ߵ���J��X�᷑��y�d���i7J�J"�8r�(A�e%z�� �t�t��c��dq!&�BͅQ3��������Q���YIcU��|�H����e�Rc�ӗ�'n;*�/�G��Γa��k��-�:VV�/]����)�$���������j�c(�j{�z�g[?�_XX�������I�ˍ����,\^6�I��{]�U����h�d�3�%A���U+����c.���k�%�����^#�̗L��]
X:%P/�u�G�?\�ݵn{]K���s�c��{̲φ�E���.�����;X(�Z:D�=��3��I�L�r��]ԥ��Pߛh��ҔV.y��q�:���ڭt[
i?�
�W~v�; n��)ϫj�%�ĉ���I���$/�5�'������n����m�F{��POBuu�Yk|� Ql������W��Q���i����t�c�H�F�J��;��$K�!�"�EJ��妛[ x�ё#X�Xg�b����Ԕ��qx_��V�"������K�SҰ���F$=j�qY�NfQ����� ��8-��;��[0�-�l��,�R��̲L�@��>j�R���c?*mQ���#p�߯AϞ0��H\Y�k���_4=0�@t
�z�M�px��^y:Qux'�La���{�8Tj#�\D9B�耹�98�l��q([	�~������c
��FEk�~�Bc�^9���>��i�,� u�}�����A��ô�Z�q�{
9@�fB�+�b�-{��n��`2�?�K��S^����H�9�	��`�]@$�p��p�T��t[�$�Q2[�٩�`�B��
m�#�t}�<��/��o�5�X����a�s)?�i�
����g���2{�i��zT?���08����d��y-�ԋG���@.���u��,sG�a�G�������V���:~�1������X����e`��<��	���@3��R�յr �y/��y�XHb"QeE��� �0�rG�$�ϭv���Y�|`������TfNw�r'����,��G��Ρ���MW2Rr�����G�u��l_����j1���e�Z��T]����t>z^T�0Tqh^T[�3))	#Y�H:w�W�A���Lɯ_���E�������#^�X������ⲥ��Cs��7�`����$�/q���غ+���Y�qε�J�,ĺ��q0;N��y���`�� �}��S/�`�K��U)��+�i�׭��l�9��5EO�d����W�<�{�zu��n'���A�Ļ��]�I>���>�ʵ��"w���B��b�o	ah)�YAhKM�H�PV��u"����"2rl�vC��X�w	��/���qh(��ȓO!!8���sAt�za9V�I�!�i��6����Nua=۩gy�~������'�ڞ1�,��X���1$���!��uo6Ԛ�b֭E��y��҆Vل�at(���朣Sj�;ZFE�{M��.%�H�<i��{�S��<R�ؔM��]q��\�E�\ta�_B�/�\�-O:�F�-\^��kYzU�[lI� �7|-�iZ����RdT�4j����	ͯzyU��J^)� L#+SSZ�����\I�Ѡ�^���ia�/9'+k��?*��xsr�9_��H.��x6/� C�g	9߇�Hc�8i�� F&3�}\˳��2���t��ȋX���l�d�I��e��ȝ�-����PH>;�nf8`�M��M�eΜ|���?��`8^۴�Q�Ӕ�CH� ���p��I�����v�����E���eSy��us'�	lfp�ɣ����y2G��J���_�����6�FF�
v��Sሂb� ���am�4�V�Ы��C#��^,��D2�]�A�<,��&��x:Τ_^�a�k��]�4����\�2���ܴ�Y��?��o8:��04�������*?|^�Ѻ��:e�,�,���r ���T_@D!��,@�G%����]6AB�3`c�ZO-�#08��,:�#������c�T�.����Z<���s��kC����֥PCi U��-�^�;�B��b�����e�ٸ�'�Q����]��6[��Q��,ź����6d�W�3F�T]���]���ְ��̏��6*N�fT��5H�
~�Y�[��W�L�\��
"&�b&`�v���^^�o4���(��߿�u��907�����W�(������
�ngg��6�c߿pL+�NN��-;�6K�J.b�eK�>'��G߮���o�u��[��^���6�=+�������<�^|)���j?�N��9D��a��-��������zi�1xy�d�Gɱ��Q��lV��ٖ����ؚ�~y�z�P�9����Pd���Cd�k��W��l��T�K�8�x�m�&�9�p���A;��*^��,��ҲX�$���>Ȅz8�0�ٖ2-e��RA�A��]+c�5ȥ����$y�L�iK���(X3��L�(>�`�h����~���)y��EEE�Ke�*i���+"22��v2�ttV�2�q<Uw�k�U��X9�{W��C���5�$���Jt��s�c��梯;4�c�.�����仜w��J��~[o�2�Rf�~|i���u�{�4�-���U��q�w�{֟��h��(4B�T��0TA��^)�k0�};��]��3���y��C,��m�삂�t%J\��m|���Rmm�֏�]�fݪ4��پ�(T���5���YR���ln7/_�s��y:
��*&X�\��j&�HF!��+�؜�r��`(���ϩ:\��ٝS��C%�y.+.�U�m����.��Q��A�/C�c���D���ySc7�s{�KW���!����ŏ!�ێ��N]{O��t p��zF�B�H>��3�׾a���m���;a'f�yď��X���1G�r�ix(Ǒb�$�����Fm'�S�U�\���&��WWÇ�z]'�~��Bk��|�)���p8���c�A��;��y����������ߟ���:7ȱ=x��wc��;J�0��q6/��QX�f�.���U�L�y^�7+$e;2��G�[@Eټq�4H� ���tw(H7H�K�tHwK�"�t�"�"���]�����Ι{8gٝ�����uϘɶ�E���\{�}�7�4Y���o�o�;�9��]���Gy� �B��ɭ�i�� p:	�G��Ղ��L	]�csu����MM�"�����\��^�Wb0���Ƨ)�Z�P��|g��x��o�F�9�,V�ڑ�����{��ԯ|��S<��orF{����A�+��^���SMM��S:B��)��px�M�*X���Z�TdR�����I8�kR�rL$�'j:��U+K��e�d|�}{��2,i��÷o�*�5�x򦿫6y���:\��uQ%��=��OÆ�5��]O]�����T++�U������]������UW��zZ��B ��ϗ����"c����Zb��ML�0��⣣�_��LxR�O���в�7e)�����r;$�Ǌ&�����i�2=+>֞:9;������#Z���  \�d��'�n�����u+�����N����G)����������z�����P�u{�<e�9�Q���NMܼn�R��m+M��M��a���"n�z��x��Fa��F,ӂ�����D��M���#�Oƪ�E>�F9����4�j��Q&�u�Tk&�ͫئ����T�N���Vk=Ѱ_RR�jP³L<L�ə�"={�E �K�{�"0a�=���n�5`�LMԎ}����2=�~��@F���x ��\ӵ׵�w��ATE��� �%�Fֈ{�B)�?W*;���K�V���/�6��M����SN.ZԿ(t֦�L��]�E8s�[�iH����]b{�kH2:
�m$��I�foZUJ�h�Ij���G3����K��M5�Q��yٲ� �Ju��e4[���",#J�x���vc1{@�6�ʜܲ� �;���-��{f�-R¥�[/�L�]d����|���[�:����02�Ҥ߼W�r~��[����U f�
1z����F_�֫!�=J�-=!G��u����Ϻ&�	ϯ���TÉ��'��!OW[���}p�A� ��	䲠�M����c\B��ť�����a��z�7�3�[qC�/�D��R(�x�:�$s����tx�Ջ}�(d�B��d���q���8���ʭe�������u�v]]lS�m&7<���W@I5ߟ��W�'��Σz(z<eR-�|����)��\�<��������������ޮ(o���[�)u���cqy{�����=t���l��9$0����5��WR��3G~S���Ho�{�LpK�b��Ȩ:z�~9cE����*���ɿU��Ըc�Z����7SJs�_�GӢ6��n,�O��!�N#�ɘ�.�!�e��?[4$���9;]����M!x��~��X�Os��`�5F>�Kz��'�e�^Ђ�Tc����x���Oy���mf�S�2��ܟԒ�����3�4@�Gɱ[�$f���ϒ��ۂ
��"��[-\	���\�~Ϯx�R][����o_�� +r���1��_���*;��la����{Gr#[�Q"�����vѥ��h6�����#|w���"'ǲW��,������ �Xd�V&&�kڟ>�e*�V��������K��J��XM�yg�ۨ|������B�Q����Յ����~WW�f�x��/R�gL�lYF�X���'�'E�p=�*�W>c���fs�{�&#?��$Q��N�Z~嫝���N����k�֐︕z����T�8LhV˲a��]�_
k%�vB�Uz��
:���,p+7J|sx��t�� �ַ�1/�sǽP���sU��������[��O�j��_I���]a��=Le}�gN�?L�T+RCdrg�y�������_��Ԓ�H����VT(�
�E�ک���lq� 	1���ַ���w]t�V�!E���p���8d�~���������Q�:�<�l�����enn���"U���z�!:&f��[Hy9��V�X���d��(((t@��c�~�����p7��a%��Z�MS8ꦭ���z��H���:4�imS���W�o@��0�}�qwuq�N��O��	*���i�
X��+a�	�1C�.f�3�,����?��ba��L�]��T�z^�Z�����"*� p�{j*��@��T�5><�Z�0��q�( �
��^�}�����w��4��-n[������xDRo�\���|��*S��L� �9<��e�X��s֢Y#G2�]"�R����f�k�z��ב6�Z�Q^P��I����װg<c(E<��f� ���]�����f�8�k{�B5��>�j_��vfQ�@u �,L�a�'Kv/R���p���q�HYۮ���ͥ0����7�ګ���LݎV|�{�;T*99�x
���i>�!s��H%�~(��iJ�/<k�V�e����MX��.r9���G����֮D�_��͵��+m���A��&��k7�M�벏�B�� �ʣȷ��DO�{�U��	n�׎�ɝ�l�ií5��,~|Vũp���ם$�����������[WL���_k���L͵[��O[l5�2�Gs܊�����S*@\v��ŴQ�D��Q9��,]ڈ�F�����xȥ���K�l�Ҩ�����G8�1:?~`o�w2<�?�{��W���N�ͶKۑ��N�Q�1��7�3't��^S0�Y�
��[��-��ބ����"��f����i�QJa>�h��P���I����v1gљťҵ�G��1�����?<E���$x��}N�-dn��'Уۻ煌�m�~��?����΀��u�~�������l�h���K,��`X}.&!E}Gd|�Z22���O�>w��#�Sg�Oj��l�Tppu\/��^���\�q|�z�^�$j��sI�O8��ށ�Nv�tb�<�O+�u�6�+�.���>���?�lM�\vJT0���Kl��mg<%yS�TaV���w���@���ˁ�ҵpip�; �?owkhY�bf��kh���N�Rl`)Y�i*����eo~^���GŌ� ��E^,�UU-�Ga�ށH��%��t�b#���U�����{#Y+I>�֤]ta%�T���9�tr#���3e�D���Z~C`3X^ET����a��F�:���� ���zd7<����6���ԛa*m��k�|�Uz�Ӽӂ�|!�A������YvwZ$�uw��L�C��yC�ի���k2���=��i��m�͙t��3��;K7#�N:[,MC\�؇\�d�j��/Hd�>.T��^���f��Ȩb``���������0`�c���@`=�>^V��y>�-�\0�-�)ɲ�I0��9��$-$��ejxz�_�����w;�c1aG:l�zT�?�����-?����S�S�xΩ�Kn�(����y}�¼�:��{�gHhf���:&�
|J�釣,�FN���CL�ﶆƇ��*R��nw�۪���r��]�BԊ1�2���A��?�*uO_��L�_�2���a��lU�ҟݒ;���k��u~�ʪ��a��ɗO�Ƌ��(Q("��_��n�H�P���lL0���,rA@�8�2�P�7ӰcN�RM&
k���.w��Jc5b �Յi0�K��v�e��0y��"z�ud�8͇��>�]e8��T���=�;obf�$�R7x����c;EMd�C�q�T�v�Hz�,��X���p�ZׂR�����)C�n����բ�֬3�j���Y�w��^���T�l���'w�t�����ǵ쯇j(e~{��im��+���@h��/3T�IIH��z�"N��U�9'�KS7Q�Z8�<�^�
�յٳG�|Zy�f�4��z���!�s�`�w=b;E�-���?�8J���������kz�д��[��A������piH}�t�3~������	��5>O�^u:O��]�Fx���U��$b�,3YJ�,�_��[:�ߣ��ݮ���R�k�A
�ܭ�eCp^8	}N�������MMX�Iz?a<	mK����+�-�t�r�%I$P��2q��ڡ^af��$1��L9$�K�N�5 �9U�VeU�m��O<�����o��a�
P9ac��{�~`"U�R署��0!h~qR"��#�~����V�.S�\�r����b����O��%1�@�oUUx���"W��U �,��=GG	j��yk�qMމQ��9E��k$3--�?��{	�E�h���i��$G���� =Y�)sp�}�H�����x�]���K9���q$�߽�����GO��M��JkR~b�}���i���t� �V��̘%���?��6$>�D��6�������j�� r؟y�� 2�#�*"P�9���G��v+��B��؇Ł OU��(����N���c�Z��*����P,�="_>>�f�;�8^K�?���]&2���0���NQZDo�z�N}4z|���;��$�j]�S��~Z�MO~o�j��q=�Š%e�.v�X���0��~������,#�.i�/�*]rK�Y�Zy�G��}=��cf�7�o���А��4*<�c�1^�d� ��wq�k�����+ה�qg�Z^�YQZc
p�'�d�
�hQ����ػ mˆ@fj,qΙ�7/<i��-E9G�:�c�?�)��÷�a:ޘN�١�\��g���=h��f�قV
�>ڃx�h;|n�S+XlA�M�qT�M�����ݑ��W���i��18p�Ә���͘j�[z���e�?�|�cy��j��Q�uj����WF����ă�@�,0���&���S1-�Ϻ��{���a�O�����!�h9ҿ�Z)��ـ'*�����4dv���k���h	��x�e�Ǚv�n��n=2&������A��f-���~[�\���d����?�[�߄�#fe�R�������-h;Ƚ�o��/A���"��~p'L �fL��&�H���@����gv�*����CP��/ם��>/8tam�7gZs��	猦ډg2}�R�@����/����p��(1lj���}�Դ�F�Wh�M�P?�Xy296j�!;6�h�A����U�n�Ջc�FG����|�wf����5Ͷ�ca��n�>.҄^������7�6���Է��Än���j��]�FM�6�X�:Ժ�s�A�Q#zBBC��
�`Q��D�jX��[8�kM*++� ������P ���W�lZNEOxB���(�Q	��;�t7�sR�2k.�Ӯ폂܊\�35�A�[]i\���5�~ch�J�h��̠��D;GqѨ��A�N�Nw�c�zSPh��d]�t��O�Oǹ+VX�m�>�����a�铻/
��؄�?��B�H�3^5s���q+,zW�a.cڤ�]�>�Ƙ�n�鹈�H��tQ�O�7Ci\�|�.�IIIK�zqey鳙V���ҸHh&��V��@"���愤�������N<��5���ɒ�'�o��f�@CB &&���I� _�;�Ķ�嬤�X�2vG�/���E���3y��.[ޗ��/�ڒ���,:�S����`>\�,e�~��aa�l�X�~%��Ĳ�H���ܮ�=��vz�N�VVV������K�g�ܼ��>D N-δ/]�)�zcK�z|5�$�G-jdL�����H�e_���E��#|h:<��O�:��Z&����j[��[��8^����E����,�Ê��[Ea8lW����k1�X��h�󛶥�M^�[���#��:�g�Z/����7���޴�Tk>-��������T�>�r���}�%�_�\�Ч��r�LI�_=>>ZS��������c���28�g�Ib�Ј�Z����\�����,�����v6o��L��bF�d�Fv����j̜�k"O���z��q���Y��@"#o<����C��yy��{{M���KQ��^���{	3��m^�f6�$�u�*O�ﾚ�(���o�g�T��M@�s� �E�������8g`�݊_tz��R7���J��OJ�+���a�9�������U�&��ƭo�h"�Hj\�94���"�هP�X�#��^TTG���:;]Q\�������$��J-i�W���݋P*��{p =`�T���gu�������~t��:�7��Gz<�NB���cY�.����w�rvWlEֶ��Tf�lw���J����~+-!e�sVl\�FĔ��M��z�Lm%]����^�YLU�%�e�e)@!!�.�lV���9�]`��+���y�y�j��_��=j�뽠���e���xx�E��|�y��x�������j�K�����$�,���"���O�v(k2���ۈӈt����<|�r�� ƺ��B�2��G~,��|�v4���$�0oߎ%��)�!{��_%@G�w��(p)�5�H>�����O�~��U�����:ɿ����؃�8�bw��R��]�=Q@�N�?��S�J{_�%,�{�yOƫ$ؐkK"\R.y��R�x�6O��>�.t�H%�5d�ϡQ=�ss��%�><iu�}����YJ�����`��r�y��O�tJ$�v�r��8�,���6�WȠ��w[�6�7��6������#:�`q]`�ND3��e SWͶM/�W�h"x�U��$ �n0]�����������+g7��/J���j�"��>0��pĽx��ɋ�`���0K\\ ��Hj�����'4����|�g��ʚ~rlaJrQob�		)eOA[��xvd͐^������6�6�O^k_$Z���-jv�ʹ%�4lĴ`�5�{���?��tMeEK�PD>=f����c�<��2` ��8c�r��'�.'���#g)�����Y����F)ܱ�&t^��]��0څ�)	��b34}����.����gb����`�P�/��D�����7n����P�@I����Ns���e�؇u��W��\cI�~3d/�����Z-D���@�¼X��T�#��#YB��?�Kh��.p����nE�f�M�"R~�-��P�Yt�)*�[G��:�R~�	-���[#A~u����̜�6�:�����T~�$);w��p춠��X�˪�I�TK�9������g�qW)�{�K^�%QϮzc�)����w�Oʘ�$	���	�q��桡ܸ��^DˎON+f�v��޿K0��*V?	��ڞ�.:�2����:Rs�:,�,����B�3P�]iiSS��n�ᦽ1�J%��u�z:��N��퍕��R�?L�=�_D�+��a��~�zS����KR1{:���[ڴJ�y�9���BD�pp��%^ԑ���Ͷ�����!7��l�x�t7A������?��ц_��L���(���%��-����������lU;:����7�BJM����hU��޵cOh# \ �|Ê��w��'��Q��Nҁ�KYB�i��a�^���fl_�����^BCC*VG���� ?��E��T����B9�M��]��~J�������{�n�bu��f#����Z��o��|�t��$x��왽=�m9>U'�Ѿ^�j��4-�U�����^����nl��<�U��rd���.�}V�Wy���&9k���K�+K����Q��&�'�����gK�?n�q����@$x�a�g��?h�������qI7+B�J*�Gk��>�E��<Z���F���.B7�$�9p[�X�v�	?��^�Q�򥣴n��G\��Y��;T�6Cć	�kS�Vچt�A���L�K���G� �kC=y�Ҕ�&�#^��KI!��9o<髠�Ɍ}4�]��7n62�Y��~��2S���n�y./|� �1`ط"&܍b~�7�i��D���c���%�����e�غ8?/�9����<S�t�R�j!e��'�#�
ITS�L݉��Z^�I�S�'�7��Ȼ��"I��5�
�ف��E'j���u��c�	c�t�����&�ol�� �@N#c��LB\3T��|����D�����A�(�7l�x1�յ�2�f��Nh���ZP�^�5�U-�ʞ����y�k�*;B���NGS�
�Ю1W��h}6�i�i�ơ��6t@X�>�Up`e;Uک��	�F�N�[1l�O��O�l�{b��;�tB荈�gr���}?��Ղ�K��):k��4��E����O��b�",�s�)<Ї��^!d���=�Y�P�c�v�)E�.�q�Q�>�]�������jJ?0�3�+I�Z˽�I-Y���ngx�@���g�"��dW�Q��5(n���A�o�d��(C��_/�Og�dg"#�Ƅ4��<�i<�ͥ��j�Z��	�Hq[�ϊƻ�]!D&���d'9�����e{�مմS<�e���<i���ߠs������D߼��_8�>w�49�����gU�-�L+���F����<I�Tǧ��@�y������Y�A��,�~�^����M�vf~n����z��-�w|C�˽M
yG�ߍW�`���8��C��gf~kߝ�ZeA@����
+PV!��O�q�_��ު>�u��X���g:�����y]ϚB��D���-.t;g"�-���!bf��m:N�B�j�mצ���L���Y���5]�n�'�8ł
�g��f�gp>>>ڵV���ŏ?�kL��y ��G<���cD��Di�s��*�Ol�ZԯO�,)Ը6Q�U{W*	���)��`��*;�s0��W.<���aV-((p��ۻ��7_#[/q9�Y3�YH�SaJc����Y�怨X:��)i�
�Ɔ��>�pL��ts=��sJ��gCv���j"��({ݻ�~h��{�}iHqsy�>������nV��~��+��{T�a_̆�x�JӮf�_���,�}!�)�R�h�7H��V�6�7#�<PX�kC.d���[JV"i�*�~�☥-d�R�oޠ�X���(�u�,[� Mb�JH�ݽarcH^Q�G�7y�S��;�Ʉ���g>�$��r�)�+�|"�1�3e����(?��Y�{�??�I��[��F�r4�; u`���A�0p�F�&�fJ�l�6 �g���u��~�mO{�Qa�S��D�~���]t�cZ��c���I<�w�@�nP�����+NrZc>�nP����r�=�x��I�=��j=�u�xSY�;���>�X<*� &B�p�y��.�Vр��7I��&����8��(Q}� ���v����t ��:��h��N� ���(��I�bfA#��j�'7�P���N��D�[ ���� C�y�q�Ix�Ȑ�xJnR>! �śڳ�ꌿL/�I{o�p{�в���e���0�v���Ne���1$��*��)�^w�N_�Rs7�E��>��o85:���~?T�ڿ�S"���ykDFK+u�\噖���J�O	������5��u|D��W����@W�|����~S+�V�_M��?�i���R]�;z�\�^��N�^�q�K"��r�tΧ����	��lX�їH�]�{���L��@�7��w���nݳL+��l|>�*d><,*�}ቶ`ta�����[C��I<�w	���5Xc<���<�_�%F-sm�-P����% �8��p�;yR��`�j>��Ɯ6O��8�j<�f	q�A���ay!��E�9�e����PM-1w+?I��������s�Ol�Զ�/�m���{<��P��O��	q�H����;Us^^���+M[�R�?�_ӜN��V�;��m8����f��ַ�1�ϓ���~}*|r>�O:dZY�~Hܘ>>2͟��5G^��v��#9��Ϛ������'��$�Ԙ�,JG-�m�a�~�^�����2�݃e�as4gPL�5)�bҷu�*ޢ�m�����>CF�s�ξ�
N:�qQ�n5����-��`K�b�	�r(����	�Ҕ��t���"���7�&�7~#��a֎i��*SX%���� 5]d�F�9Z��v���D�?�9����Dx%�����gw��f�R��2`�\�О�B��Iǎ���H{wtE�7l��^@�n}�S���������LK^�ʝ��)����P����䙻��8m�F!%Y�����0����eՍ�U���\�?^���F�YQR�kK���q�A�H���d@g�z��z�H�h�h:1FI3G�+X����
t�h{6�b�F�����sw{t�+Xhd�v�Ш�}�p�+��UڥV�}��z�ۂ�o1���ʥ�B�{�U�4�G��95釸](1$��w�Ì<g�]��nI����b��f���f���p�mX���F$Ϳ`Sy�����t[�p�40dM���J�E"��Wz	E������\�o�Nə�g,>Sd:y)�(���VO�b~��{��Phx㘀�T=�v%\�fُ������͝�5)<�Ir��+薴����!]CP(􅺔�+ŉ�`*{oO4	(���]�P6́F������u.8�����F9��/zȀ��g����p5�l�&����pɪ�%��4d�>lUP���,�w��<�|��Gr��b@:���\�ݑ��Q*��}��@��ޙ�m��9�;
�<����\�k��W�<���iZ+�ʦF���cLI5=ފM��N��=�<�Uo
n�K~\�H|MQ���P'��x)�؞�QyC����,�ט����w�������c���<iJk8�X�K.�[q��O����*𽈎��JU��m�,9���˻�>�byY�0�N��	-�3�����|��cV,T4�{���n���Л�خU��Վx:�8��J�n���ZmM�g��V����|�~^�2��ꯊ�����W.�A"�aq��q"43�eq����}b��zk�Ǭ�߯�����A����Wwm�#�1u�N��>�㋓�y�k�_��|�[~�-�9p��'���mA������Kt�lE����)h����S��V�Z=�^7�Ӡ!S�������TŒl_x�24f�L��\}�� .�#'�%4�dI�/8���d��@|/Xu��gl]ڽ"���Ɖ���;��p���s��R-�J����&�缾�wS�
W��e6J�������=�w����hk�?S�*�k�]�Z2�pK������-�ul8����Ƌs���{��T�t]������o��Z�긚�'�����,�i
Ps�e�.b�doN�m��SZ5�d�O�0��%�!�>��eR�dlv����mB������M�qL�ܿ�,�7</���Лp�}�N���8�\,z~t���e��yߚ�4G6^�"�[�'�ָF n���hk
9͎R�~'�����Ŷ�u��%�������)M �����d��-�\jqS����T���+R6�&Yn��1����L�l�}l�
�l������ߘ��������>�.�o��Ã�}uxx
p�v{����`;���%qKZb�����e�@�;�R鶾�>n8 P�ʻ8�����D��m�//I�X �* q���o']�٥x�|���B�
 �H�ɗ���X�6����e}��]�3˰'��Ӗ��ΩBE8�F�_�(�M�ce�U9��#�����7�'S��ˏ(.|l|(c.ge�e�Pl:/�4�2���xb�K&]1ݥh���{%�����Em}Ո��}3�RlZp�J|*����Cii==�͡����zG�˔�����L��a^�;i�^�8zy�OO�.-�_]�>�[��~��̽��H�@���(��U��mԠ8.���~�g��-�;g�=�W���9�]�-��:j�h�I����m� #���c?��nK�\�N��<�'l4���ID������ܒ�b[��!�1}n�ٕ\��	8��n	�>���\��lo�,��A���E������� ڧ֖�^5��9�������OQ���}á�%����c3r�x�U�In���s[Qz�w0Y}q�碴Y�����/|4��������R،�h4�=@�a�n����U,�h�ۏ�����~[j����2x�F�Tvn�M�v��D{��"����DK�AC|8YYY���?�S���?�˞)¬�f�@`���^ 1����S�mlG$����)�>�(�F�W/�>
�[V%��@����h�s!��ᇯ��'�a$G,6�Q\Xh��aśhN���"adD$Q���N��3U޾UJZ��Z�,��R`{�V�^^N�@��������;;׬��abaFcac�.y'�h5�L���c���:bu�c�Mx�����~�IC;K�r[t9�J���(`��+�S��@��i���skc��Fv���}g�~�JD�u�%���'��F����.5-Ĳ�KLCy�u3[*�'	v�x"k'd��%Q�jӠ4�j��O�q��
f_�[f��D8d�?b�3u��\1�Qn���$�r��Fy�}w�i�(���8���y��D�'�\� �\���\J|�L		�g�T��:Y[��	u�A�����斖*�Uɡ1*����&�b��Oo��]:�,�����擲���L'H���EP�"�ot�5#=�����Ԩ�׎0�0$��dQ��ȓ��<W������x\ny�8l�&�hdv+����Dc�r�e�
��L:���5:����yyd���	�b�������q�<�A	A��o�G:�W�2�d4E^�7p�ʴ�nT������٥c;/����"��]54��ꁎ�/��/h\�%�s�����?�W?0�i�U���	�0��8Գ�34~Ƚ�� $f�?����c_��V\��Ǎ��N������ �f[�L����m�6)e�����]&گ ���-u�dK�.����_,������Y�칏�-������T�f~@�K�-���c��%x�f�!�e�<+C-�6Sc�u��)U��t9�t��4����[g7����\�Uh�]ͬ]����k�^�}o�gsqw�ki!�k !;�:���ׁmԄ�P����[��7�ayUUx��O�����&�zc�|����I��ǘ[}m'ݩ��6jt���^:V�4�T� ��0�3��ݧ�u�`��\�h����.MSkA�T" 
�)26��(R��ǈpC("-*�3h����ՙ��l�iqѴ�5.2����s>˷��X�#3��@#N�%I�dJD�+���� �U �>���Y5F�A�SaZ%�h�;D���0��Z�Q�K9u?�k(���ʨ�f��P}v��Q�	k�|�6�������#Z��ؗ�^_���0�����c�F��D�u���xzT�ً����$y�"���7����vU��MNjLaOB ������W�����h�ՙ5�E3�Q
'��v��"-�K�w�ĆS��(`D�'����W`Wm �:�H�,�;�``��Zo.���,K���\�di�d���r � ~�C�nB��nF�sss�l�$�P
8T�Ȟ�,�X���Ԅ��8�K6��Ⱦ6S4����Xu n~�O��rl~rl��?�"'':i�Q��l3�\9g~��+�:XX��0(=\�`�K�q���M�� ^�1}�Z\��
fӄ�P��S�B�.��=���U�8I֒n�r�ґYBo��N��=@e&���i�{.8�Dm��抰E<bF�(���=���䁋n;�Y��-��ba�τ�b�"�h`���w��Ld��֎�F�����-z��l�R�B��I��d�
�Pd���s�ZA!����p={(!���r����ZG �L�=�/�3�7��!!(,��h�J���{�B���ʯ�¤�	�Z/�΅��&O�+g	v��(�w|j*��vJ�@~���J�&�'���FO�n��R���i=�Ȃc���<�iŶ�r��E��� �(\S�R�].���|$�\�����Z�x`>�����E�n	��~�!�d4��|Ohu󇍡&�}�?K�Yf�`ۃR�����	�z�˼ܛu�I&�K�?^~��s�Y{��hmuZ]u�d��VV���C�H�Bn�`*4���¸�D��A� )d-�=��6Q���)<�YK���$��n�YuS����))�1Wg븑��c�L�_kve#�D�Wf�i�g5�p*�˓&j��R��X;.���	߫*[7${k�ٻ4�����2=&��m މ�o'+�&&�v��v�N�u.�qs���ꇣ]�V����0���e��=��b�5���VVLG�4�DsB!���2hUR���ӈ������542_l��������1��l��7�@���R�+�����ʸHܼ��/"����lmaxP�VbӨφ$��h2 c�Ud.��!�?�~�!���78��+KK����1'}�������Ss�S�p7��k`���`)�k�J�;h�(�j�G�x�e����e�X�P�����ѯb��@8��~�0��nBX�$�f���L����O:�m��8�r�$���c*/���o�\#��m�NJ��ֲ�
�������W�·��=Ӝ��1n,DRc2��� �������5d8Ӥ�I��O�вx�	~�!�f`��*�����(��B�P����J�QJr��`#)������|U�Ю����g_Q�*���0��H^{<F ��^��5��f�D,)Np��Ԡ�a����n��W���ë�G�N�P��qݒ�S#�[a-M�J�,��Q��<�v-�O��L1��yv�TXe;��
@-���$��n�*�@���0���`OP��(�/�%��}���F{e��7Y����kҗ�4h���d�8Q�7�����R�����Gc4�υ&ma�\���o�����q���\&X���
�'iӈC��:,,������"�{z�����L�+ƿg�݇�o��L!�~Ǝw����>�4���%ڏ�	-�Iǀ+oQ�˔��#���������&�ca�4y��t���;�?�W~�����?[��u�߹����*����)����̓[�wFp�ӿ��j��=�qT�I�E���k�Y^t%�T�-
�(2���+ݚ��+�f�C���Xx���,����vx�W��Ayzo��O� �%���چ���\����#&R���"�m܁�K;W����]}�9_j>�O���i����
�to�!�:T����IZp�_ǎ߆++6,8�}�;����=�����g�n�#i�}�4�"i!d��|=R���(0��'��TI-q�xؼ�0���Q�z�d.�+�|��c�H��T��!�"êj���#;���W��A^:���e��-��zΙ�	4��i�HII�-��N���8��mf�ˊ��f�xU�?�0z\!2�'�[	x/������{>}r勲6����t�r�{�EFEB�Ks�󬐨�~z� �z�Y�W�ŀ��m?1>nkkK0�J��[��;��Ǯv �Z[�&o�,1-G�5kd��ǋ�{�skn-�p�:O��f׽��m>O�2�~����N���l�=N�4^Aޫo���&	@T�qBP5��`�Oa��0�/Mv�9W���}��>�шh���>��F�!	!���������s�aBP�at̪��ls�e�O���2=�[z�7�T���q�N��Q{�� P�}n��bH$��n9M�ǔ�[L �ۻ;���������7G�/�z/��b�*�)���a݃�W�
��߼�	�O�>m��ue[�C���3���Y�����]\�m��x_0���r�ָ�5�I�,�)bK��0~]"�e�~��5��׿�Ѵf޳�ߋb� �AB����)¢a�W�|(		�]!���t��3�+7�U�!�� Y�.°����S���BjZ��(�7 ��v`Z���V�?I�w��'I��ֈ�=�/�v��K��Gb0�[4�F���t�p%N�kM=t�p̫��Z	\���A��E � >�
z�3����˴R�����&oA*�ccp�X�lw����CU�i
�\i��v��) �=�O��F��19�ϕj�\N��nM�Q��t��|���z��Z آ/�)N~`���J�{l�ɡ����畦�3s��?�|���.�A����-��4��X�Ҧ���v����3�J�a���EM���8���8I+�g��Y��^��N�C]�	���ThJp7�"�\:H��	�ѷ�WU�����w���!��(&&�d�Z��ٹ��˅(�H�܍	�Tcb�I���O
�l�aE�Q�*ue�t��_�X������:z�Zo��m����/�yB�o�I\J����!ʰJ��֒AjYD�����~	܏�`
���Uߐ�Bi�R�&|�6
�"�~׭ؠZ�[�ȧyu[�7��ء[˪� ��L7,S�)�!Lq�,hh�f<�*��.��� ��m6�p��#�D���n��Q9����H0��G��I]LZEZN��fD��8�͖���S�v#�in,�׼��c�@|��a�oĵ�.�kNjf��ΰ�v�А�����l�|^_���u�������ea/�|d_z�̮�*�chW�>���133���o����xc3l�
ņ������͘�e�Y�@��o�yf(��.W�����ʆ�m���j���/��.'p~��[�+��B��L��%�\3z�-�r~�(S���&M7E��[��|�B��?�3����,�����7G���^dN�/}c�3f��Z03���}��u�����v�q3x?��԰�Y�YY0���ͤj&J� ;�2֒�l�p
��Vvv�^vV�!f��)��.���@�<՞y�20 b7��$Z�ʹ��]r[r�[|�#���<�-F���҆�o^4n�Ko��u\��������6�&Y��D��j�J��l�ֶ|ww�֣�Az�*�?����M)<v��g�'��d�}����[D&�F>^^p]!@�o�Л��I�ߺ�� ���%�NK�;׬��E	! ܲWm���
�*����/ݍ" �)� ��"��Ҡ(H]����D��A���;/���1w�q_߻g���ٳg��5�T�g{݈�ϟ��:�Z(��jU�T���)��߂��WJA�0먉83'��'�Odv��u�~���-_V����Q��ܙ3U?�xy�[�
��k7�������!�5���f����Xy����I'E<�WW۽𶴆���G�A��1WWY9��gm�h�:t�����.�"hRFٿs�����ď�f����s�v��)gc�B~�5�eH/��p� �'œ���� z3^��
�h1';��;n=|K!�J���Z��ݧ�5����1�o�S�f��{Wҁ��	a�Q��6��p��m��HM�S]9%%��SV�c��Ʃ�#�h�����z��)�̬���X��q*.�<O�<��������
�a,�0�3�t_�[?�X_j֛��5�g�����K�k��qO44K��$��NE�П��-u�_�D!��[��$�'w��=F��;Ư�F���A�՘ ��	g�IZX�}{֕�ض�� Ha^��X1müX�z}����7s�X3�'O��0��t�^V2���T���MR�O4@�zA����i-�U2������_�9��v�z_s4���Z�^W�	a� ��,.�zJ�Ȼ�)xT��,�J#g(!� � 5��db�>@����, D9I�����O:[��.�n.j.�����*-�uRw��X��p$~��i��$�n����������t��i����	�����.�
Y{�Z~�`k������R�=#����� �ڭ��|�?�1�`����;}�d��St��̳Z$;��t��唜-�����]e:��Ч��ӓ�����[�P1��&�PE�f\Q�e~�l�H����3>�a]e�F$�|�Gq!�y���Ne��bD�j�8�l�$�hW#7:�Gm��Pބ���̵'L/t=�)��;g���>t�})�c�]��E�6"qCΫs�U��ϯ���ï�ő�Y-	�Ǐ>�),��p3����.���ֺ�/}+�!Ұp���B]��x=`	�f�e�	���B�i0��ˀU��9�6_0�v�fg����ؽ�2�VR�-�?�s���i���T��v�}�����Ϳ�B��``���D)�yA��<,_������M�Kꥎ�5�J���=��W�Ax����&�XyKA�qn�o����#��D��j��A�t�j�Yy��c����|��$i�ae�G�� �� ��� t�V~0é�1��tL�'z��H-�F��Uu���΍���~�aאˌ)�Z�+�=��w�ҡuv�qa�]�~ w�7����4�]��V��U�}�I(k�F�����}�uT� �D���=�����ā��^F�3�����8���[��E���Ʊ��tHt�O�~7
^M�!��� ����h�u!�h��P_��:nM�����v��E�W���H`xG�쩻hף�1z�����YYL��+$:X1�t�#+�!]4�g��}[h@��V�g	�h�-֏4�X��z��y��L�PU,!!��֙DPx��
 ���E�Ǻ����!�NNvwS,���?��P�X��-�ڕ~����є�� �[��qzͤ݁�����A@9M)i3�o+��.%%�K8����Bw���ȁdӂm-tJ�)��P]�ǀ��F���Y�	��_�)!G��\�a�-����9k$�zQP�I����@X�`,I�3�w�F<tz����bɨ�QS��Q�\j�ܼ��hR��n~#�p�	Ob�>Q��^��	;�S�0K�S䖎9r��X"!%�뿋��������Puk����`Dp�1�����m��F�4���,?��޻
S�w|�M�`�p�-De��b����%`�^^b`Q|[��O�3��{޹s�t��3�*��B8/����a������&�&rҪ�|M�.�{������,�GB�/���-��<�Ѫn9���5l� �gff���S-�8tj^�\�|��v�!��i�G��ܐ7a�����p�ef��L)�՗�$E�gϰ�u��mz�� '����SL1I0�M�G՟Ϭ#�����b����G^�$��uQn���fswFj�f`����lƉq\��1�Je�̸�]m�i����8�0�F(t����H�љM��1�5u��IW���#�{�fo�O����p���#��Wl���x�1T7�l{``�Ǵ��Bk��o�tf0�i.��`~  ��>h����6��*r��U}��QXXx:�"�]{�z�q�_��՞k�sa���2�����/����@�� !3�L��p{��f-+���D�Z<�]#��jr�y�驩�2/i�;LL�D;�57�/�m#�h�Sa�KHL�]֑�2w�/�� ����Z\��I�W�7ݰ�hӟ��~�*H���8�OɿA�hP_��k|����g,�N�)U�MI�ە��*ܛ96��/��B��d������%TU���W��uՅ��ST
aď�)aI4p
Y���v�߂��9Q�i�#�+6=�V�:`K�;a!�?׳ޗO��no[Ae����i�	�6����ĝ��&��������M_P�V\���n��yyy��}K����D�}�~�����P��{��^@#h�l&�������;廉�E�pݫ��`׮J-,�]�5'h1�(VI{�2�ూU��#f�3a���S}�Q�tl(mc�f���`MS"�>�~5�e=�@Ks���=����j���KQR�A�uW��4ך�R�n�{�=9$O�|soϋh}Ua�ޏlBe������99������#��4>Y���z�L�������%��)�eE����9�iшl$̒�'mW��|��̡tW���\�2�t��ns{Z^����٥��k���Oũ�{��\�Ə��L�h��r�?3Ĺc�Ԅ%/���`�F��= �4��r�x��t�H#�U�H7B;��̺=ڮY�(�=PM���L��>����Ђ^I���|�ߒ�a�3�A����ڵ@G�W���К��z�E��׵���;:K|��~i���d��E���b��ۭ���*S^}�Z0�������guRRXS'k.cc���8�z}� k�%����v(�ڍ2�d���&��m�e��P�R�vq[3�N��ԋ3�3!��8u5�É�6�4��n� z�}G�a֒��yc1_.nJ�V��C�o"�S���7f;�ӧ�\�5�4L	������A&g�~Ρ��*����Z�ٜ�Zu��+\4��b�Nc�F������ޙ�|�����R�1�3sԤ��1K�1E��+֊�����C�w.΄c,}G�9jJ��(qN�ւ`TUS[�u�i����T������[�#����0:�!(ck[�7��<cy�з�̯��N��qOO�徔��i�գ��K��$,�=	�����ә� �Gߣ�q2h��R�6�HÝ|�/�/�,�a w=���H�A���;m�|�#$K.æQB�����0��"��#�;�Շ�_~��I�h�R�|��̋>�"&Ts���'��̣@�F��\�[��a�[��冕Z����.�8͵��R	���:�6�J����frC8���P�~��Q��ɘӴ׹;L��>�b�s����feϗ袕$�����w�׼��x���Hf���ˉϷMJ%y�"'\�X2�^�B��
���{�Z	6t�A�>c�\�3W{���+r2�GnU�,##��6���f�;/QQYٲ�r^^8�6 �SSF���Z20�e�������}�L����'Q�ݙ���r�:�k���<�������-��~���JK3�ѭ����E^���GL�^���+k�$��i;��a� �Ԋ
8S��1�K~����n�%�+����[��s�-�]���d}�F?����hi����\YW7<4�I5�KLl��o�A3 �%��q_Y�P2K6��h�'Fk�l�{�dl��� &����秈�?l���mL��;�]?��2���4�J�Hܩ��A�cu�p���������I�Eo�+T�s�-���%���\}�cag�1�}$dt;*����V���)|4���˚��2�b��-޸�8$�c�b��<y�o��+��Q���B��F�k�w�m�<��T�O�>u���P��5�#''�����@�ʊ���@��p�Ǧ]�F�9Da0OGIG7�G�]�G�f���bDf���g@������5ϲ��[�4v�&?<	�Y<k��g(�u���MXF3et���W<����%�����>)|����Lã��]g�����T̰��8]�t�T��\�	%e�b�G��V��P�E�M�@ Jn�.a���w.�{�4'yS�AB������W�K�?�ؕ�R]ܾ�x��r���8HF�g����IX���g��W�N
��e^��)Q�lQr�����k��c��CS�6?ڴ���U�+B���E.je.R�M'9���^@�F1��l��`z
!��8�oLL��z8�V�qӆ��^��� ����CJJ�2���UV^�707	���+�������*���G�{����%44ځ1>ٞq�-�?>N���wQ�U��>~oX���Q���c�I��?������喝��I�QjԞ�B�0j�Ǐ`�8����K�t�ӊ�����~f�� �e������qK ����|��|r���?D��O��Th�[��b"ʔԬ���˽���y��L�d�wOr02���eB����3S�L]����Hj��˻:�����Ҍa��%���6�S�5p��X��D��ê�5�K��F욋��B�&��'g�S���J����'T�����{�Ԭ�b�)��o��
B��b{S5�2ql�gi),�Q-,���P��[Mr{������b���+yy>�ԑ��ߑ�W3cE!h������)A���eM�{�C��B�p	�A����^A��w96Y�Ⱦ87�k?�]w#4-*1]]�>�E|�JC���So~���{�^����Z= t��L��<�'���Y��ﴏϿի���(�\J����,�L�U�9������?T�K
)�C^�`M��Ϧ ;J(á����5?�r��yXo�7!d�!**T���%�'�LHv�Z�d�sՇ��Ž���3�C+OB���	4oL�����g����3��uW��̹���?Ny�z>�LO'��M~�.:xN�U�H�M�1�N��'�Z|�s�ovl��o�"�χ��$�%x-i-5#�f�'r�'�$�b��������o�����oGJRDB^��àr!`�SũV�'k��ЙŪ��3����x�4�Z�-X7���({��)�`+�`�Z���N��K��E�K��ǚ��(�*!5�e�D��xQy]m��c���䊖~<j�CG'x/|��E�����˴ՙު��!����G����5��O{����Ѵ
�>��~����%����s�.�����̃_i��jz���l�)Nc>����s_�F�NH �:4����+��P3230<�!`�!�Od(V�*W��oGݶ���(HeKJ����6ڟ�zV��&OJ���0���m��z�-.����g4���ǎ����i+�[ ���H��Қ�|(�Ց��.4V�:>.n>����5 ��H����y��l��	KYGG�0�ƻ�l��>���X|usSآf�QZ��_@@���3���p�Y�Ռ��~=��r����t�Ջpi��W)�a�N��ncsLa�"�p!���uH5�K>��z,��������C���,����M�s�����%�c:U�nB/~x��~_"Ǥ��N��h��+���ȠF���r�~�jH0$+���@q��YW,��{��*�lS�P[�K�g̊��PH�7�[�!������~7Կ��ύOB�,����*�������	4��v�JD��d���~`fF�[�Ck��r��y�$�ֵ:�����S[ɇv?��ao߽�NN���'�hUw�'�'�?;;���G�����F>�}7��hhh i��-[����	5�=�3 �F�6���>�#,,�9	���v�L��A���J�(����1g���F��:a5j��?�����(/��B�&����r!&J�
��y�wNJ<.�k������e�o�������h.U�uJ���wK�8,-8�?������	 W���MM���y��Ӭ�R�ڴ�۷o�'&\��̡ҵ�������CWLL̗zz����k.���Ձ���\	u��Ӄ#�>��M�G�{g}^�I�!������G����Ñ��S�y�z~q� ��ۑ��S��,�%���=_���1���fN]��kw!ܯCƨ޼�|v�F�-��o	���5�v/�_ݵ���V���)�ac�����5{N���a��m����v:�L{J5�Dw2|\ѧ�%�*��Ü��CThT�^ ���`��D1���U�1X�O���^U�|����f�[p�`�qd�P��xx)���T��>zU���K���h|��knβ��b ���\�ؐRT�-x�&Ku���/�ܥ��-���N��7H��I7[�h3����n�j4y6$��� ����`���m��r�ׯ��� ��S+	ߓ'�Ӱ�]'�8�<���@
�@>Q�_�A����G.����jU>Q⸥�ܠ�9^z�G��#�ѽz�
>�S�x �4�;?�������b�w{�n�U1}xN�V����	��a�K�;@�N���72��DB�8��G���d��%[��e�
�T���@�]]Ǧ�y��8 : Βn�����Ӹ`@x��GD�:'��GD@��:�����FFƚ��B{�MW8J�g��>���o0����1�]�_�᥊��c����lM`�N�
���Q����M^�w �O��"'(*++��QQ���M�Z�Գ�$?�=�z?a�I�ug;���I"?��3��r"����#Wh��G	`��y�����t=\���dddP��)^]9�y����_�9ƪyg���?K�m=����?�%�=��E��(_opV�3x��G�ϭW:�C�u<��|=��| ���z*���J>�ɛAH,�{LZ����eT�>[�����w��9�����B�°�y�t�[�4�������6E߂�YV�>r�sJߋfm�h��� �ST����B	���]NE�+�/�-%��^Wb���;0G������̌�R_�i����Xm.���j��ni?)	w;�c�����<G��pa�|N^����yI%%��+�	�,�%S[�VN�Ɛ���=�2r32��yB��Rϝ$T���f����aI�����eH$��j�:>z�]N��Bֶ%-OCغðУ�]��g]D��1}BBN5����}\|<�w�GiلeHJVV<	]��w� ~�VU����;��zs���|���,�<��Qutա��R�K�D���%�j/z��=��W/6�AE�oM�w�	b9 ��O'	)�4b����$��F�j�/�R3R�O��ÖԞ�f��v=w����\�M�uc�8��H��LHϴt4�/Rbo�쬞�DZ��N�O9��_(��$�t����N�5y�Gc+���e�'���҉�ЂBN��$)�p�\���`�x��m]Z,hck�=M*���m�a���3*%O~��1A���t����P,|�Y8��PF[�dYi��-�»�w �K|�g!�+3�A�%g8(D�FqS�8M��Z4������||�Ư怣�R�RTn�� o�5����MM}���X�y_�֟��^�-�H�锁�x?o'ۭU��������߿�Vd ק��ze��� Rκn�����>�U��[aҤ y�/�Qe���Ҩu焎�P��ǹ��L4�ė�'jpF�މ��x�M��q��h��tu�/v��s0w�� N��EP|=��S��SY���C��Q�-��||�E*���j��a��0��Hˍ6K�PIE�RRZ�G
P �972_&��ѡ!��9O�<��3w�$�/6ˡ���O�i"���������d��Lq#�\9��b(s ��+�� 3#���X:��7yrtl:@d*�72��P%>Y�s�c��!�n|�̸����4_#5��4�U�+��=Y��.M�g$�]Ao�4�&��_��0!�ƦC䚢�>.x���>P���9��D����Ϥa�;����ϳ����O=A*Ey�E�6��Q@JrtHߗ����4C®��Xg�W����}�m�w�5̫� /+�7d�0����KE~��_�wL���	 9JO/g?�����sW~
\�7o���[�����cs2��(�$�p~��K�?^.�ZקK%� �� X�2��
��S�z#
�ѓ3�����	��v��GO�M��Ձ���S�˛C�եS
}�97&���J�{5nR���W��W=��hW�bs�Omv.)WR��v��w���A�V����B\\6ߐOV���*���e���>��&h�;�����S�s6�i�вN��L!]S��@hj���'#W�Ѐ�r��q�?6�B�'���RF�ݠ&�e�ѭ���Ӕ���=���U��v�ٍ��qq ����ޡ��&��/���F{=,;�[[%�]V�N/W��R����]��7�g��TS�v��;s�c�TΚ���n��P8`yM^7�8'�������W'sr�h��J�?H�4a��eU��Ed0�(k�ZW0PQ��jDի�*�
s��:��-�9��2��5��}l�f�@�huk+i�I��u|��J��I��xER���T�JI�̎�F	1ƕZ���r�ʴ�ܡĮUi����G ���#i{V���>Fď�_��1�{���m�8]]�Uh���s�֛!&�����:��89���YB�~����x�ص@\��N�		h�NkQʘ����� |����8���OU�`��M���W�k�k��.� ,�U����ee1Y~ol�*��7���6��FKZ�P����բ0֏t��O�g�pT�����(�ƀ��.�	�ĪP+�)E��U<[��9��m��<�k���kg�1�q�vS^I�r-���3��DSP[QsSٞԨ����XF�#��)�y��G���Ma���ש�4����BG����%egg_��	�t����fE���*�C�� k��SS����or.�{�5�|���8���?q095e��Dk���x]�m����*P]]]�[Z~;>KOO���?��	��y�/J�C-��[�1g�󡶝8U�`��e'I�4E��(I��}]�.kЪ����Oq�c���������g���܄�,'|��%���2�3<�}#��a��R_���I�e�n��8]0܊���ö����4�F����!��tK\�0p�c�$���;�6{�VqRRR ��3p+��!��aV����7���x%�ܾ//T�֠��l9����������DI�ﾗ��P�h�D��U~0��	�CiN���>�Ϟ��7R�#�G�q�#(�
-@��6���%�_o�Xw��w#@#�ۭ#�� �&�ߜ��ӧ�8O9e(N\ӫ_l�l�{�I�JL�	
����>B)�{�ȟ%UB�Sttt�L�&x�%�G�w���X����^���Ĥ%���Hg?��V]B�^(�SB�"�u[�P�4(	_&��q��m���y�'�4�|�٨u=K(T���qk1�W�WTW����l�t����*�Y>Q �.�C�UH$##���${�ZXI���n���v xП�g���L�d�����D�r�MοVF����KW����fT:?m�0c%�wCy] �RYYY&*l�R���;�f���#1���̟�]�ޗƱ�h��-�|�{j��x'z�����2|�ݏ��Xh���-d��_�Bxe�(�p��L
8���������;��ܗ��C���fD����k�
4?C�K��Im��`������ ������>-Ï��f��#X��#��#Lp��_[�� �9ӢJ4��� %lQ-�MY����lmm�Y7�%�m[ �CH�P�'����p�\O��7�8��A����=J��vz=v�ڀ��Qn�\M)��';r�$�BY,��Y̴��c/�eM{u=��r*S���/w%�x��?����'�x7hK�n�>�2c:���������a�γ��%�ł{�V���(����GAW;�}��̛��)��?#��g$Q�Q�|n�n1`�~�z�P|ͽ�vR��,�%y���4dd�:�y�}f�D��x�_����ujE������ �ml��s(F3܃�]�H�'�U��Eb������@���ݷ�2<�������2�t���i`��7b��jj6�d �]hb��8?o��uT9�2�7k1���"�$ l��E���4��A�\ �^&���g��_3"���?NA��q�6q.��]R$l�Ψԁf���1�0{v��^��<�صC:���$��E����u$7,�DB*�ŕ�S-
V�)���q���\�*JJJs+����Ϧ5:��%a1�YO��m,S�*c	��8�G
�&'S��_T�����!$�H�L��q���%��	�N�GB����p)���O��̀S�^U�HH����v-j�VvW�w��V�-��N��q�����*���<��O�4�i����ލ���e6">Y���3>����,�_}�6��i=;�7��o���e��t͢'M�qy8�2�Kmq�ts�Q|+���,��o��]��9���������`E	��)S�������A���f8X��&i��w�Xo+Y88 a������2)t�	���iz�z"
h���J�8݋&NB���� �>��Ihkk�XY���s�zG�o�o؞e��n�G���p�$䴸�N0�w�9�<��A��������l�T'��)L	�I�*k�����T�h1�l~���|�E7��ۭ��vE�kb��x���Nݦ-`���(�\Z����ص�Z�"*<͇�J%Q��لݗe߇B��a���Y�>44)B$6��0|\G.�0�R;ne�}i杚.(]���"z��Nf��5]r!�Bۢ�.�:��z u(����5�K��w^y��mU��N6�no{6Q�.�455���	_>��[���N��
U��4ݡ��ݠ���[r?�W�w�HGO�P6��~����X�n2Y��.뗗���T���a�.A�w0�CT��o��ıoQ�����e=�0x�����L��G�P�
Oۖ1�m��� 
:�A��EB� )D��0��ChBƱ���}?鿿o�#����6V��{�i�@0���_cY&� YH�"�������B=r(���;)����/�L�gb�zY7�� ���@�=�(N��D��d	Yل-�能=O��f��DW��_
0�Nǭɀ�m��s�W�,��,/M��ܙ_�B�����JV���1%�d�K����NNN�Bs�)�j�MTFR��ߣy����UWΣ"H�+���=�Mj�W�Qiؕ���|}���)-��ʂWՠ.���^�F��i�]�H�;	�3nkg�� 5b��EH�A�\��V�K?��H۵�H��v�~��q��?R��O��ښO�A��׹�����CUi�8�
�Λ��4����t�tCɛ������r)i���L��H�{�� o�|\q��?���~R��鋤��1������ mP/�H�T"��- G?5.g����q/෬��o � �7�!���%`�?�|�ص ;09�h����0�r�4-ㇶ\�M��IRz���Wl��I�?o�p�k�Cϗ�ME5��K�6��%��}�'??ߦ���ْ��"\�2 ��ޝ��&���t>]�ߦ)b������	���8w�]!*�@��Z�E)Z�equjG��0c>Z��%�C#��O£����B;Һ�3�{P�V�Jr[JU5́o�_�=�����Z��Tl�Eڃ'���*q�"+��pqe�{�F6z��{�Ώ6lk�����=�Q�����k����Vb�MǕ�A��̣e��E��M��2��W�,h�A�Wz���"o��������r����r19�R���
#�#��F�$���)4��vb��wE��1-G��*"*%g;�$Š����¯�Y����MW[:�ܨ�>�Z��9;m׮,f%Z�tq ��0y�:�ˋ}�����y��O��ƉaRT{֋��I��To�o�V/٧9�nF|����;����B�8�����x882	�����v([|Ѡ� c=QĽ��'�CK:���i�9?%�y廯�$�D�7%l��W��l�JH���|��J��8�	��@��x�C�;�<�>l��H�,-�^�k&j�����s0ʷ>���/���9���eb��U�(4�쥈o��a}+m}b����K�0�t��쭈ݐ�"�3�+,�sq���@v)����ާԠ;c�:��d��4H3}�D�Py�K~���ǒ �%j@�FR9�oN���7�F���COA�&�˗���n�~Q���ݘggg�mi��0+�zL4�,I������T�6��ۻ�U�[4�"k�/lY<�^��Yu_����hQX�SS �xr���%���%�D�F�mPJ�-Y}y�e�o�p����)�P<c�	Vub�ٴm{NQ�uA�)�;�-!8�@�8:��p�$��%6�R��A�~�����4a�"�p%�=�KO1�[�_^�ʃ�j�����9̞ˑ�䃽Nj㡬 �B��o����Es��v���,�$�������<|ͨ���r�Ho7>���3�Ϧ_z�st���ix�����Bs~q�	�S����5q+���3I�?��.��N�8�F#��Y>�v�.���ܗ�Ӣ�/��R�����1�E��Z �'�
�{T%���_���g� �U��w^��` � A�-Qd���1��/^VV6�L�TE�>��!��Nyp����c~~����;�>}z�*/-�sbf�S��$#�f/c����h�#��y׀�5�d	dt���7�����"���!X����.W�m�M�,�:�S�tg�z{:eȒa�{�=�^�v���2��Jwm��0�����X}�BA4��b"�F!�-�İx�
͇Vڳ��h$7X�Z�H��$����	
_�n)А��iEii�������fO>�����A�2B���kH�22 ж���8!��2�^(/�����5؈��<���r��z�\!&�]����<�*N�@5L5���[ �}�,�o�p�ma�p�糿�mDy/2���!�4����h'��k�����M��Ԧ�����!cQ�L���O|�$F;�1��"��Ux�Ɩv�B�c�@!�ЁZ����q���CY����s�Y�Cj9���Él:(�O��ѾM��e��&�������#���#��b���_���E�^��i_A)���.R�o��eNi�Pt�G<�aۖ��&+�XX���������^3) �L4_�)�)���#yj����!PDh؜�y!����>����Iv�R�Y���������g7w}Ij���[�=j�K�$%%e�E0�,�f=��:���񢍇"���w�Q��X}iXj�oj��NXL7� ;��X�p��f��k��7=���]�v(>��Y�Z���%������G��߭���Sp"	���ug5,�W��?m5�h�;C]d���<���ք4����|j~�^�5
<�qV
@�p�\#jIn�#/�o�H�cf0ڛC2��� Z�ߓ�	����U0���_�G�y��O��|��;�'nН�� ���6#bB�2�>�3���X>fw�]1tGV�)阮�h�f��Lh7W�vN���J������7�bUU����PQ������3����]�¯�=����ɩ�iN�����ᖌ_=w��ώz�"x�s�|H�VK���,>lły[�:>>��y4�����@�Aw��2��*�4��Iw��<̂��]=�,�9��{	�Y�w��{F.ݟ�4����`2qz�8���03������ʶ$X�b	z��:9R�_z@0�:!���������J��ŉ�j(	뺩�R̝s�C	|e)�h�~��pR(��İO�|���Y[[�΅��{�	��4�`t�����*�(�AU#*�K�n��������@����%��uP�|6�.��pVm)�ՠ��t�(x���h�\O3IĐ�e(9��C�L�ٳ����zL4��7��2I�l]E�嘛������y�|�.��\��A`�;�'g?n�����&�_����I�S$�̘������H�?j>��ʧ��HJJ2\=�g�a
Y搈��ʍ�MmS^7�J�����\���1o�"a�#y}�_�	2�_6�/#����E�[�?�.� V�����[I��`	eaa�p����ϛ����m�[�y�!��x|Z� 5���9[�X��:�,�?���3٠)��u�N�Z��\�T����2b A�����#���O���",�ۯ}�"�囤ǈY�jϏa�-�����͑<BQ�+m��O�	����9�#��2��Z���Ge��RC��Ň��O�	a��P�hG����vM''>��5GU�@��4�=qorZ�}������F�Gng��9N(��x������^���ǭIJ`��g�T1���[x ��t�R]8�"^<���n����w��Z����32���
���,|}�U�99BoǠ�.Cu_�kA#�IU�����qG,u����Wz�j�>&���*n�>?��s?�'3NK�^�K�R�tlӻ@��GH.=Е�I�&e�*-K��vz�=$�W�LO�M��WWb�y���b�-�)̈�B�=//Z?������I�m�$��` xi�P�oKvdm��t���	��qFH8�Uhݑ^и�Q��>����-��L%2�ĳp��´��N��]׆��⠹���b9�N���/��W;^�"n��I�Q�"BD��5�@'u^�* E�c^��ί&�É����h�z4l��m"��B����x��\JA�5�78XV�Vs���!�(�� $]j�NN:}Z%N������#�@�)'�����K+��|ݙ�����$x����������H�͜�}��oi����i�>�>R�����1���z?�(�>}Z��"�]]��뭭[D��L����@N���`��;�(������y�Ɔ�\+��.��2/v�T��BѤ�zT�O���fW�ݬ9fㄵ��v���0�D��3����qd�<P�o�݂U���L(�ʔ��*c�Ujg�z���v>$3�}30>��<4��O|Τ��9G�{DUU�`k�� �U|����p]]]åc��qi�n?ړ�8�[��qk�g$7��(��o��j1���>E\�ɿ	w����F2j�4�����m��3�
|�ۀ��"$��UҜ�|�HN�G;1��]�Md�����r냗��quS�������A�����?�z�/�W��5f@�ˁt'�x���t��"�0^�Ǳ&LGGG��ot�9������gr0�5�5;${�!�t9�˰)�&9�0�\%a42?»�w[;.no�D���ɹ�@GX�����ι�vk@��B��F5'08�ő�V����u�۲� ���B���PVx�[JY�?�s��'Wb�1�S�y'�e:96��ը��Ą��fƬ<��Y+��(&1t���]���CE���v���C�U(����ȝ跸o\��7�\����-/]�m��F����,�e���r�hp�Q�Д���;�e���}QN^?��5�@8�L�@gNȱ�}���l��eu+�2ʰ���{��.������n8 ��88-+��I���Όv�l�+9Е�ʖ��$��<� �d��0�$ۖ��c�S������h�[�y�H�vY9�S@�����N����k)�u011�fB��7�}�n���-b�zq@�z�d�k�~�^X�߆��{���3���H������%Y��]��F��[�K���fq�������%�KP2���E\����e1�f|+�E��Z���j���P��-�ׅ�������hDD(�I�1��@��a�3Zl�K����hd��-}F��'>���"f��(2j#�L�&�50�������œ�_�GHGY.�C~��}_���h�8,�+���N����^�#��P�YZ#��,�д�R�3�v�X{�N�q�?��:����^RS
�;r%����o��wN������h�M����7��_;ȗq�^��j�V����mya�`a���!C����Vj&@�fJ��\\\�O�˦�Cc� ��-��{vo�+��~w*�K9 ��v�۟��(�W���%��.�O%�dY����50@��C��E&�qq&!�A��=��gԮ�y[�8��AFQ�]�����	U�����60m�k(|4�b�G�����A�A<��r�X�/�j^�1��IH'^�C�O�z?c�,c�^"��cMF��,�j��)lQ��z?@�b|s}�a�͎T�� �m�)g8Lb�,���n��:vr�(�}�{����ô�,��G�"\\\�	O��
������L[��'� yi�K�A��@�?���6g�%b�x
��vw�m��\�㋧��bL���ݾ����8���0�	�ݽ�t�賷�3K���-88�#PeKFCC���A�Y��k���r5`sW2r��!%%�Z�����3u�Z�D|��w01[�^���}���v�NU��s�g��x�#T�;=��x��Atuue��58:�I�]=�H.
�-�W�E5u1�Kn�S�d����I���}���9���k���[�P�ޤ��>��t���ߕ���⿚���gb/v]�a��b��yh1`P�Y�^ ��T��ⶈ�-����ϊ�K��oZ�=�aZ��L��^V�e�Dz�/..ʷm	 ��j��m+�J�.Z���]_��+ t���Zz�|��ML^�y�|os�3�����,w��승��e���o���z�#����E�b|Ǆ�������Q�XG�`�7f��Wh�ubY���	X�3�4��;�O���g��pH5و�-�r�b�`����Ս��vR����>H����N�A8}_�aT�L>�'��SS�]Q��a����)�!4�VY!����y���!���ܴaY���]��Nn]]�ZF�fЗ,������7�]>Q`�	�<D�+;}~�İ�P(���N%y�5 �n'�@����d��})�x�]7
kNf�J?�5�^׾�~�Gמ�����9�x�S��T��o�]�l���d|w�^�$��*|&fy��tϞvQ~��1�PQm�ߣ^E�t��tHK��tw��t34("�)0�t� -94�1H����^���b����y�{�s�y}2�Z�ms�^0w4AHL�QUE���՚Wwl���P^^~�H-�r	�:D�R�@��|%N��� *�C���mS�����A�� ,�w��c2m�g�����N7o������ò���,�X����- �km8�y]�k�������gO�hi�#`[\���"b�7h럳y퍾��黗����-���+]]�]��m��M���{�j�����C�}+[��SY�Ι��Ϝ���?Zc,�y{X���޾x�S�Ë
�h�9U�n]��A�>�DVYYh�,��:w��=%���߿�G�0�@rlb��Ϳ�����5 gNc���������B�s�{{���(Y�����C1���!�9�A ��ɉK����^�5�Jo��#SS͓�o�i����P�1sy/+/���!bz�k�؊�/ݽ�}���+�Fl��:Ek@*���� J�}�*��$�mU��K{'��cQ�֢���P���.���&�i_�� �_g�4S
�X����8�����p�{6�^D�N�1<,,������T9�o�z��r����(����<���$���RUK�ᡡw��$��`C�J3�)��cJ�	H	ş6������f���'�H+���ΐ^^��rnT9�����".>����uyhwy#��5�'�[������E����_[X|���{�Uo�����b<��%�ՙ��O����:�i?>^�M3eѭ�!b}�P¾����nn�Y��L{���"�GR��4.�M���⟒�ƽ�IL7�n�EQ6,��UD���Zj��t���-����6==�ck���{P�۾��9Q;nF�	�l�k�P�qXO�N����TM�>0�:��Qu��!�����E�L�-����V�2���/�k>,�3�$�H�Y�����~���5/��ޞzn�{^<*����K���č�T_��s���b��5vx&hY�>B�t�+.�|q�V��M�vf����;�/�У�*�f¶&+iXYoC�\�����W�`�>�>�j�ƠH����L�i[]Rj�`�h��/Dd�G���'{�!���jñk�^�ץ�ͪ����;MF�.���i�RDf[*��(1�9�y��5)YY�������w�c�0G���`�۪�JRű�4�di_�t�	�c�&�֍���ަϦ_�2���X-c�ڵ��B�[�����}H��?0?"d#{���<��t���5�l��e:Il+�X��bt?��ܨ���^��Ds�L������)^W�c�_'���w���ձ�����m���J�û�%[:����+��'��̳���c�j�O}}E+lQ
t+��8��{��ʐJ��q�څ"�3��Уe/0gs{=���Vo�AbzM���'�A�7�����a^އ��R5ؠ�c��+���}��Y܅@�Ԕ^YEŋ�gK��!	�A ����nQ�n�xi|��8FT��F�_7	��L8��c��J��/x�}�d6�]&q�ٿU�|�u��U�@��b�M��BBcbbn���`����ҧgV8�(|�{��_�������>�.��Շ�����GBz{��j*O��F/�]�	�����������wo���ߡ�ލ��`O�DebbY
����*ъ������{s@��u�w�+�����;�僟��?Re���	^�q�q�|����e]���|��[���~,��IE��0���E�]S,���=22%MM���S�8�L[s[Ҋ�_(����.�����J���I����l��O�b�AmI()%TU�ǣX�@{ʐB�~�����z,229�7�u(��~�0(�le~&2侥p��!���5�k*/�$+�o*"?"���]!�	���WRQy�������@����?�L������z P��*r�Yŝ���T`0��m���bq�����̎�:���~q1�@+3�5������'�i���@�*')D�Bw����
J���n�m�����-�Px�py|�X�\d�;]!�$x���'C?�����b�p��5f2�D�b"�#�tX��]����e|�b�����pZ�f�(���T������0���3L�g�]�����a����ar�����Y�x�3Ӣ��ܰ�_O���qG��mZZ���p2�cE��U�U���Ó�r���	C_x�P�=RH��&6�R~��i�Y�:��ۯ�A$��~�9P,)H����L��k���]I��^��'5�	=�������X D6�x��s�Ҟ%��D:�ë)B��$$$�/T��-F��#�L�4R�!����Ѽ�������|5�)��}����1S�K��h>�/��H�����:d|��f�b>83�x�����̬��F:4��� ��P��Ʀ�� ���۫пTWk�џ��"��!2��t{�Q��J�b����?�9=�j��p�-��6KO�b��):�[��>z����N�	�Q���)?^1ʔ���XGd�KRWQy(�)���g�a`�ê�EnW��(r��*}F2)�`f1U0�4 �Px�i��[6�3m/��K��� t?�>Ya��E|��qq`�MMLXY�)���
��o���J�_�;iJR��ϋ��@h뛛jpxeMm���t!��iQ]]]uC�"��Ng��?8�rf�7�����unO�zɮ�WM�2��=��^"�N!�bd�|����k5��d�<�
I�6�IG��R�?��{�}]_��;Z���c5.V�
X�(D�����?��σ��l):�2�&T=ڪ� B��:!͈��щ�i�f���ɂ�\&W��^����{�]K��t0#��/2N��}�V�L||��r_��əut��
>S��n�1R@Df��%�0hV�1�?π���P�vS`����I�����3�Dyee��W�u3�܏|��f��[��Z�܀ݻۡЩ�D��z��icfb�Ty��q��9?~)�ٽq`���P��uī�_�|7�lϫ���q륳Z�9)���ۈP��3���o%m���h�iqj3R��Άݵ ���� |�����$+@��g8�Q���U�\����c��Qwy���Ht�{}�6H����=�Тmt��n{ز�P(�.�����	����\Κ/x�W����}��|���S�U/w�,��n5�Â�<2g�RI�w� ��ڢ��Q�����,����S���8��Xuʠ^�u�R16� �P�3o=Q��=rM;y�����%�s�s^h���h۞bim��\i��.;XP9�+B����%$$�^�����R�F�����bx������Q�� ��>����Us7��g�=���Ū�k
�D�����1.�'�Jj�SO�����y%�tU2j�;t9�t1FT��y��,���50��
Li�_����*�N�\dOT�V�U����Qt,7�7_d�󩇷����̶:;ܒ^�_��355�̼��������Q�����z�B"�����`xw�j�����8����쬈>E���.A�5����-:::��_��M�lUL���L��dq���	� �4u����N���>��� ��,��2 �QN}§E���!�Wa0�w$ab���V��=��L3����պ(��!}O�t2��|�B�z/�K�C�L����e�a�R��>-��3vm��Ѿ2{e���nO.��SR�r��!O�A�����bG�KQ>��2�x^�x<j���p&�,�n|�%v��5��~������1�7`�[0V0�d��?���������p�ә�m_g��$���A��q}�O�!��JJ�G=�{���F��0�tv�|u����E�g�k=|3e�t0�{��ޏ��N��x��/j��'�t0��'����EF��2>�%�3"���,�����$,�FX�7���JlW�����C��kF&iPV���ѽ��ֺ��Tac�}}o倴('G�ǧ!��i���#  ���V�o)�>�.�8N	 ��v)^")��8��ibAC@��	�E�;�a��O����q.��v�Aäʒe�sJ�d	���%���\�?�����8xr�.�]������B�3��p��j��{��-(Pם����ܗ��8X�L�m���C����Fn�֎�f\]�Eտ�Ю�����D�7�:�(�v=v�d�F~uS�~�_�A���#��uk��1M��L�n�:����u��c���[���܁$=
��;/[�c�n���a9Zk�iu>?v���yd�B�f[��4r�����OH(Z�Z�0s����w-/m�K��T��fi��g��B���k-��j����� 3���h=�VB�w�d$�П��/'^�M�IMY�ܛ����A ���y��+w`�!������1��|v^�l-��X�|ζN��Rٽ�d?��[���8"ǧ���<cI�O.�8hZʾ�O�����������8�S�?q2KI��x����fPV]C#(�������8�㜳+����t�e�v��K3J
���̽�~��4���4�IP����*I,�<��~�t5з�BT6�����=���@���V����Z��ޓ�1�ꇋ|�y_��j\��#���a��È~`"+l���$--=�{�ʽޠ@��y1����g�pD����?Ж�vSqʙ�V"�����>[B3*Η[Z�ǳĞ�0_."�ˏZ��HCӲN�Ҽ�@<��B�B�eD06:��lZ&��Hx�ǽ��
.3���aԢ�	�5� U��!1fă=��AR��E�S'�d�`j�����F���{p�����~��f��s��M��mo�m }�f_�߳ �Zk*/J�b�ު����?گ��[�S�����dt�K��r<��5�`�&IRRr�jtC��˴�N�Ѿ��~����v���~�}U�E䨺�s�H�xS�a��T�ZU^�
_x)tӻ��|T%éԹ��'U����+5q�$0�}o�b8W���E����x�S6$B=CV���L^�-��خt�:��\\\������+�i�2�HB���zD5�� ���֮��8c����%A�B�b��T"׈�q��UQh�c3ei�ങ�.0��r344�^w&����u���[-C?j�I�,���h����l�4�?�SQ_m^�K2Q�:�=����{��e�qT���,�_�S��l�:_��V�����(+ۺ>L�r#��b��(7W���jp���9�Cv�(zőhM8���!x7�M��`c��(� �[cq"��	�����[9p�/�R4A�Z��>�`cc/��`��%áU���Rpd�<��@��t�ϟr!� �¾]��槑|��5R����|�Y��3"�e[i����"r�yTJJ�z�������N���B`0�us,����g!��Mj��u<����̬����ю���d��OK+��AY���qk��`z�A\�W�9{N�����ard�i-��Vt8��n�N� {�xgAZ_PXX�˼7�s5:""M��^�v�s��KT�!.��s��}Qh=m����Eej	��-�2h��*�����:�ؕ� ��։Rs��-�,Mw	`�5�����F�b��9ԫ,y��Q��^}L��ᑑ��%.NNn�Sg���!��k���3u@5����K��4�󊺎�/,�̚b��QZ���^��;��D���oř'��Z�JUSU� s��ꏃ{M����A�ĕLp��5�M \�£Pb!�]?#���:�I�B6dע�5�l+A�������N�=#,¼��A?�U66�1�k����ׯ^����4F�t�0s�U�k�Si�TgPtq�w95��R%�*7�K��`�r�|m��`�o�*�Ǻ��4�@�� ��L��2�ܧ�a���B�Z�v"�S?Dϒ�T����_q���ZT�y�È��yy��3w����'�z0:�wO
�ԥhͲ�A��4ӟp��;���*]�׳PY��ny3j �A�DR=����2���b�V�ά�<M�e{zz�Q�"�� �.�=��	e���������y���DII	��e������xl��:�.vN�ݡ֐�9�T�Z�����r�=��ֻ,�_�f[=F[?������\K!v@d���A�/6ӝ2���,�N��H�wF����q0��Œ7C�ڴ��_P��=+�#B� ��u��Om+'A>���<v;金H�����>��|NN���p������D��X�O�<���◵>�g�P�{��Keoܓ,������ �����2�����gĒ�D�r=�y���t��f�[�ow�u �c(Һ࠮�~�u���y�=���hy٬�x>�>ܸ���Xj^Q���7R��R�(�{�vD�I���nQZL�X[1D�9�6���CJQQS[�T_�#xY�j��U�*��ط�MI8���vf�e���A�w�T���55:R�&��<�S�!��l��p^U�^ I���;B��{֠��]�'
�|��-�rt��"c��(�����I%���YY�No0/�Zit�1D!��zL~_�����[SuY\��~��o�㿠�y~�r[]_]URUU�v{����jXd�-J ����3d���üx�vi���ޏ��x/�^���Cft��}(d�����~3;�������ؖkO��'O��dD����K��9.Ɍo����᮹o�텹����&rY�=�]�5�R1��/	5]�ښ(/�����ߤ�;�tut|� �����؜��}FϪJKU=7(�Si�x �@2���C/�rS�}�vUs>\����ƕ,E
y���5�6�wȜ)����&�Y@h�yX�`.�D5�jj�����K��u�z�$����N�}���s� �0�M?wbbbz4Y9T���p�ָ5Yy4~�������Z9����65��VM��M��ܗ��l��SDX��+6��Z_=�/��ս$#��4k�^� vP����Q0�@iD��n��k�QT��H��ά��fo</��9��Kr;jٕ��v�Sm��A�4\�=�$4
c܄66�78���^���;[�~�J����\+1��2:g�ZE�l�,�� b�~ v��q�W��\Ӑ��&�O���2�'���5�F��Exb��E�Dk^�D{/7�}R8��i�ˬ�+���G�r_J����|�
��_C���G�h��(���Uy���K�%=W���A���P�[��:	��rtttL���6";n�p��5=���-��x������Q�=EB΄�5�c�2�,\`h���V|�D
��`�[񌞤d��C�I�@���@B��:n'J�	�*~��7'#ø�x��p�]mCԟ���>ꋤ(§� ���<���} {be �K�,����ͥ��O��.K.. ɏ?�$����B�x��v��})�{UZf�=����F__��):ķoJPw�nȯՐ$u�_��}��^�.Lx����#jY���U� Q�w[KA!L�*< Hs�����\}��V�h�H���3 ��%G�DH�7٧7Q�4�)3 #NI�K�FU�^	  h�nk{P�� �K�U��SPg��TPh*��g������٦5F��q4��+)��X��+>�H�prR��yfhiiY��t;0J/^����6b�j3��H���[c�'�T�Sa�ڌ�n����F2,SY;�՛�������c��G�EbAx�������E��G�	�����n�k�R�ɶ���]���;����%�W�-�ٽk� �rۿ�CFc_l)�N�c�����VJ ��|���<�8��x��X rCc��0˂IXUr���x��]�;rM}m%%�<�����i���� ��F p������Gp�4�q�����qk^��FQ4�`�9��c�t����eW�)��\���4�=��������^;��-J2��:{{G$��3�8-k�,N#��>G���.��Q�;BiM�����+Ip&��}4�5I 0,
�a�ĵ�mw�j�N�ҵVb�! �S잩���7�[��-����-d1Y��Æ�wRt�
}��D����C�QZ����~7��%��z��u�GR�j=07�zB��i�	���	��6�@{�S0�+������S
�gׁ���t�+��� ��z�����݄�ֆzѠ��j!t ��J�a/���VZ�L��o`�7�8���y�v���[A&>q�6�����v���٣3�CkDg���N&"2���aecA�d8��^�S�ˌٷ�����-�@|��0T{������`W2
t+m������j� Z����${o#��}��ؗ�YH��#G���������K����(�S̷�v�Y_2k㌝EL�#��K�z�O��#_���q��s3"���=��Q%$$��K�[+#rbl�v!���?Œ�Z��� cRR�z�R_��XbN�\�쬬TMM���h��R~C�*�'�����#�T���wD/r�C;���-�$C���LC#����T'WAWn��/u7hե�%::���켭�.�#M������Z�����Ɨ�>==>�8<t������5��,���-u�hE���M�iM���_��c^� 1��UK��v���9iii3^ �+�fD�b��u���F߯�X:�O�)����		y ����"��[!��}ް�4m{�ڤ�+��եK똾���o�n}o��p�f�rFH@���AZ 8 ��0�����WN9���6l�w�^G�e����o\��5�I�9>�S��8L�j�(��%#'g��Ǒҗ��K�s[D�7�h4O:���|+��|�Mӓ�n�R0M �V����7:�S��}�i$F�ݻ�����hsH�RO�7j�)HN���NJѴrf���
�tI��VE'�K���:�[{%�*�6	�@�#��\����tx�v����ABX�+ /� �Xn�������W��MWw7y��́���K����S�:U�i>|�2��q�vY��d �	J�١�8Q{�cg��<�^�w�`
vP"\,�\[8>���90��rn�j5��?�B�A�5'�	��VOy6쳽A�t)��K��Hŵ���ƍk�ӌ��,���?�� �G���$u���|���		�	=f.��9�U���dCkKk�lfaaaF+pi�f��O�nYO�XK)3�K~�����X��`�]�
�ݿ������N���)��vϫ��L �y�K�T�f �f1RVMI�������۫����Ѫ�/�$Z���ā�j�ۓ���(6���QI�~�۲��)l5�BHDԵ�Ki�8���q:5�2!��
�9Fn}�������Oe���{�򤴷����oa�0�M���4HĻ�D�,��J�EdgK��Q"o�M�@�6ۺ���q���=$��~�PLK����n<.F�"7��~=�5V,rF5@,0�e��茢g&�F i�%�h}h�`¯���$�L$����i���O�����g��q�pV��FY�������F�G��'l>�s��	d�ff���7a���� ������6b\�/��:) ����A�.窥ބtt��-~̒�Jl.ϖ��jq���p�)aI��ǔBnJ�L���(�]Qu���76]Ӑ�����n����0�1��5�8Ӧ�Y`��D������ţ3S����'x=_�A��BTԿ���:bV%ElF]�s#�j�5z��Hi���ϯ+��0^tI��Q		V6��2j���>�r`����m5��t*�A|?���<W�㓬Ivs�b��p�����]��)vrV2�<��u>����9����,yU��3��j�oo7M�P��
 ���5����tx�� 
�ܽ���Y���8�yu����W IݡFsQ�Yڷ^��,���3�����(d^ƕ���L�s d}s�3-��9{�Dl�'&H��!A� KOn[�:�<���2z�`D�y!G�.�ͧ�M���P�'<Y�W���Yz��ḣ"O�2�Q6@���*�,���j�m5
}e�a��􁜇R�3��Zvw��d[[5v���8n��&(*�i�ϗ��>����-(����=�Ȯ=��?+ʝ)�z��/�U�.���O0>�����������@���: 2�9dѣ�s���������>�h��s�Ky�+/&>�����}~|V��{.�Є���S��u-:�S��]7!IRe�p �>R�X�3'}�%<�m\�9���H*#UV�o+�����Ԣ
+*x����p��}/={� ;��A�\ �>��F�2�H�����/�?��׊"�I"i��R_Hb�7�'�ܻ�ڝ�p�#4J����N�cWggg�	{����e���������"Fۿ�aMW]k��F򕽽���AM^���a�{�R:�Ž�	b�Dh�IIyϊ4؅Od����X�qa��
�˃1�!Jx�����D�iP�*�"�C_��*oMU���ʦ��7�����S�!��r��$�@�A��U-����Tp}0�OcS+j��ؾ��K�����-��b�o��I�"{�}�f�;��4�H�:�ѭ���*q�G�H�9�(�8;g�?�������u+��A�o�aݟ��[�W|XF���_K�t>S�$�Q]kC��j�<�l0��~ ��;�Jߣ�T�o-�;C����� ���M&|^�����3E�!_L_����Ȭ��޵��3����� �	�F%���{�Û�t�q!���3c���*������TZ:��br>0��*$���'�5Y���~���B�$�YY��P`3i�^vE�Idu[�D��#5r��k٩bX��x艉�Wآr��c���xЫ��	 q�+��WZ�Կ m�Qy>�j���y$�&�c����i�����cia���ނ�����GAZh�=���_c��ۍ�Е��7�/Z�:�D�yc���I���E5�bW���Q����	=s5"Y�D������JVV��.�� .�0F��,��Lq� ����Q�B�F�"0�����S����7Pl�b-9`$u����^7O�uM​|��6.d�!�֮ϡ�&{!3�[*}y����N���5w.`��2i����d� ��3�Ʉ���lR�[o��H�h���0ųw�{�	B��_P "Ƅ�,%�`�,�<J���S��4P4��xI(��7��M8���:зu�2E���_�Շ%��B9�#E�#H~�k�d}��m3^"�N��"�7���v����cK���)��hI�0���u'���y�eHT�<�k�����s�@�3H;֢���JD��6X�9P�1��������Yr���T�!�ا��HP��0pX���^fg���D�o�&x���}�!�0���n:��Nni)W�4������S�w�9���2TVN۾\�>=ASU۝��$x���&(0M�4��my�8~��,��	O�(=}��8�/�5��`�����T���dh{8�#P)�.�Ϟ�>�b�60[��9%}�7^ة���f�wk�^t���o�ɭ����_xm&2�@ ���YH���T�u_*k3�c6{�"� N��9�ū�/��)L�yX]Q^��/H����)J�Q�m��d�l$4���B�o�0�����v@��X���Tl\⟝<b�|�:X� XvᛂTǡG��9�/���>J��N2QY;c��ۇF��r��մ�)H�����t���0t���Z�hYG�2�&$+���M��
�Š̑���,�zyX0�W@蔘@��
��К�j��A� � W@z�["�Z�T��ߣ=�q����{�	ч�{���{���4�7Q%*�b�IxA4�"�FF4�s�iiϊ�����rsk�}��zUL�s�IWYjV}�����$��vǰF��)��g�(�-��_��i�	-AC
�p�z�=���S�s�0ڜ�
CT�Eʞ��ѳ�8>�m�g>,!
w�X�+�ĺ,�R(H�T���K��L\\Q���U��+߾}�%1�i0f���j)�O�b/��.^vX "z��z�G��ƛ�l����ut&,����FN���@�Y_ޏK��,��KnII�Gc,�J�'U]����x����<A�x��e�篫�\��-M`���e*��D"��F@g�tttLH������`G~�y�F��L�'���^s,�������"cZ�e�ju���U%]��{��`���������:���x�h=Jg���i<I$�r�mmmh�٪�O�4گ��� ��8)ѪhI��7��Ocמ��ר5�O��uY{I�d���Sީ:Fҋ}!�EEM@o�5�9�  Y�i���J>K���S Yy�i]}��03E���^!r09�}��*\-�y-��q##�.E�F�MI���J���~�F���L6��^�aܔS�-/c?�}+�����y~���2a�qE�;�#�FU�Ⱥ��^!���?�M��F��`x]*#��K�A+9R��B�U�ooeA��\<S@%i�����.>+��h��k��Dԧ՟S�QK?{T3��2�X;g�HN��\<��^W�JSV'T�_���p��,���摁�B�!�ȏ����5�.>���qlM����#��n�_*�xSQ��p���d��W��-7Y4���~�� <Qa� m9R�xi�ie5QB=����=�t��qEQ�
�<�B o7nn�i+=�p�ǣ��{��%`U��,��ɩ�������z����99��q�̼{�i`�&�x,��%Pa9 ������)p���u��n-��w�f��Wp��o/�}� �V�,��Q!�������-RWI����q߰��p�F�%�|i�-�9����8<��o�|[q��Ϣ���*Tߓc
�}�ػjN�P)���E1̔��F���]9�E&�����O�������sO;�8��V,.�Ɵt1l��3:�K3�R����ɖۡ�7W|DAa�OV�1u��x�E_�(���f����Z�^��,��8/~
�؊�X���9�Ġ����& $�F��vAF5<ϴ������_��'_5�WiF��>l�f�R�
t���I�V��F	/ԇ!PK���E�)���^�0�����a�xL׊�[�����t۪A��[�#!~�
k*��v�������g�
����������q<Y���-t�4y�cqU����QjT���F�<���d-Z�=�Vn<�x^.��<�۷�G7���(N�q������W`^������������*�Y����Mӎnvb��K�n��\��p]&'���}�<6�w��~��b6����[��С\�)�zQr=^��i���u�)����ٓ{/[���sF�	�4��q�D�a�g�����B��h�Bo�[�����tOQM�7x�k\��?ȷ�T�r�/S�Mci���D/��O��,���TF�O��%�E=ă�h�6L���d1Ԝ����_rl�?%�G�P1�����0���|Ի.!�/���T߽���NE��rnx�L�ѓwm�*�o���G>ky��)��GK��Ѿ+��|��|h����p�BLJ���e ���b�xH~ԗT4ި�����C�a�����щ7�MD\�����Ş�3���'m��%@�dw��
�~4?;rܮ�F�R�kʊ���4��O<]�Ϲ4e�47��k+��3�{◷T�I�%�]��N Z`�Ģ��;�\�ܝ�����_'勐b�f ��Ζ���B�P�������5*2nM����Z��Ջ'�-[d�5�q�w,�w9��]5�������-�O��IU�kuH3�C�����\$9�v��t�>��oJYHL�l�"b7�N6m��G"��>�[۱ިK�w���I�,2ol�E�#���.�L�,��Z�P��&�r~�^4����T꩹O�~9E�v����hQF4	㌛�d�^����������*��Խ<[sԈ�M��n�4)c�..��{�L���h��0q�����P\+���QDQ�&��x�5�.���Y-h�� ;�m}��f5hǄŰA���R�_FV6�F����-�@������|h+h�8\���=J�q���"[b��wu�>+(�y�`jS~7������2Ʈ�b}���@iT;��ڎI���@������8�@��!?��E�lc-�����v�+�� �G��u����3����*�rrh5��Q��b�G�{FK�F ��5�=�^.4�5��v���x��p�?��يHyݷ5
���!���-i��J�Y�ᮺ�	.�X����;m�<kv��:]���`X>�i~���Fo�%���9�7����{Im�f1����پџq{�6��|��tG��X���>���e�p�w�Wm��4+�QA��F<�I��黼�u�lY#|��2�\�s4�B����CR����8�󵊟D���'���@oprr��l�������Q�F�i��uB�\��w+�S�^7+�4+T�~�UT�n-����m���zd���	�MK��*����kI���_�9;ʫK��	N�?qZJ8s�S(,���'XK\�Er�7��4p���~�ν�0����Q=��C���p����O�B���������	��l�������$Һ?�κ߳�=�dX:X?��fo��Ϫp�M'����΅Rqm?���Tg�s̟��䚴�ғ'�����3��FE�fq#O�U9�ߓfii���2�m����ѿ��t�	���#����H��߹nOD3kZ��&�4x=�������7�m��:ar�O��	��Jzq�V��.�����+�V�T���*TO.Umu'��x�k�NDZ舠auP)VfV޴�����b�tW��Ek� �m�g.��ae���B�<���;���ThƸ�:�m��K��2��~[g.k^R� ����n�̅���i�{�[�b����5kSD&qU�X]���-�X~����QY�yk���v��X�ڔXM?jŤ+�(&��L|l���.�_:yF%���f/u��ed�����i[�7`�s�$�91��}�B����Y���bA��d�4��(Ң4?��UHd��q��!=�u[��9����.AZ�i�.�
:Z��H*"kwqA �$s������<�@��%�hϹ�Ȟǖ8X�р��������tSh}�X'�1���\LVz��q/f�*������f.��v��.6�o���(ۺ|�� *6�>wZ֦�D<<�������<����"������M����b_B�(�ͽy�#A@+�����6F@$߾)����1���!L$�(q$(d�"�PV�6��h�(o�(m5Dn��p+���񝳥��n;gf��ُ�V|�GgKGg�11YO��o�ao�Zd�!%�����0���U��������ޜ��wbI�yH\�������n��dVi��>�X螃�GMJC�G]��q���s.&����b~p���@s��@M]��z�GaV}d�Y�\x���$o#��r����".kw[+o��"wX:�pW�j�L�$� �sO}�y~��օ v�=<H�`�Z�����	�\���w�j=�;�0؍R�Q6��FA8zh�5�`HU�e�m��ܪ�L��aQ:Y���ҎKr�2��ۑ�T�d�8�L#��nA���Z=����݊h�������Pf|���N(M�i�F�Wi]�g}q��Ӥ�'rΫ���Ӣ����[���C�Q����(��Nu(�|�D�$��w���S��6"���{#�fa��G�9��E� �tv�:{�H&���'��G���Q3�։���H5���Ԩ;�!m3���k��}�j{cᄅY���?<=�WٷU���5$� �m�KJ`z�=`*̸)Y����Ma����?F���G��XT
"9p�C���$�]� ٰ�ϟpb�S��%
'��7��	�_}%��'l�^^Ssk������A�xu����^;��S��'p��z��z#�W�qB���
<)uR�tø�JQ4�cwa�ɖ8m::�]�r�H��f�F�H����;��D��^��)�t&��ݲk�z.8�%�]����ؼ��~���rK��B$m�	Nf��=�)�ō��ڢ�U�~���9��G�?�h�Qn7��+٘�!֩��!fS�@�<�>���>t�&`~o�34=m���4�V� V7���Ą%�E�ʫw���fc��f�T�0*e��P��5��[��8-��"}�]�B�rt����l6 ��5�gd	�G�q_p
����=��y����(�ء�J�5>�]n��g1pc����z�<Z��i߶�Yf�F��9�.��g�Mn+�HuP������Q��~��_3�;���@F7嘑B�3��Y+'YGfv��~]��n�W�{\.lsy�y���+޴��%��)M�F;Ĝj�r3�(w�<�1�^)��w��M���k�W��}F%my�fc.�7It%�����<��3{�zz�k��Kx�ޓ�C�A��V#,�)�	�Q��Y�;��A@���J�k����EM�ՎX�r�ϒwcԘ�-�Z�@�O�zN}}���
�Fy8�ܝp<)�qqz�W)�Rʄ'��941�����=L3�j�����(�0^rv����8��,����<�Nh��:�@�><2�%|4�t������z��m%Q�75q���k������%�K�(>�i�t��6�����Z�-�I6le($�RԸlT:5`��$�y14LW3����zŊ����Jzs�!�ڭ��i�k`�4 @C�ׄ�F�q-ɼ���T������L���B'���SY�%�m��yT	_'��6v@�~2��=�f��b�j�{�_K�v�D��<�:��y�$?�A��X�6P���;S�V*�mO��u%�9;�
��K$eM �'���\�Q�Rq���8����q�[��N�R��C�^���	�er�6����씌����^љ�
SM�!�p��$�����i��g����7���su5�Lh��`�ϋNsl�`ª��*|c�rfDApˤ:O����G����':;�ٙ��qw�"+B�Er�����l`1>�D&�G?��K��ύ"f��^T��7^̳�Ч�+cm�1�����@�>��?q�u�վvsӊT30����O��c�ׯ---����i �w|��P�bb��7BP˲�佩�.�&����0@F����<,*�\*��x(s`(,�+a��{A�i��0�?#c£��feC��t�%9��� ^�U�p�����N�F����K��]�G	�Ppߘz�Pu.�=ԧ��!L�AX=��6^�b<�o��6UC0Hݣ�]7��X�M]��t��QM���^�n����[�(��n�cY����.���?���׵�BB�%CGG����ոl�JC;�S�N�+�p�ɯ�����[_U�}=���ȃ�(-(�-�"�%����AH7��0�H�Ѓ"9
�C��Đ��{/�|>��{�Aa���9k���>�И#7>j��?��.�V��=���@g��U%,����
�s�o=�l��0ඞ~Y��>'U�褨��L�:&��A&��UC����AP�ZOk�����W���g< 9`�ed�(2�2�a�;|͹�3�2kR��P�S�:X�r��Dl%`�� v��`l�&�����%���J�����rUK�I؅��y8���$n�g��<�V7Z���sO�������b�`ss�>oRhh���Ժ�q\�:���J���n�Ql���K^1�؟�V=F�+�iVr#1���ʅ.|�g:Bŗݰ�\�I+6[S)���,Ze[�@�����L��2�q�2��N��RF�?h�]��!!%����N
C
��t����j���`��� �9|i�+%��:��<�~q���̜x���]uaf�4�}��~��^�R]�~{0�E]7U�[&�cW���
�=#{�� ���S�/Ow��'���M�#��E5r��%z�m�o�7|����{J^y�}j��2";<���g!�5Ri����B�]����5�~�}�w���`�S��j�$@��5d�N\�}���u2�!���r�c.�$�M�,*��=Kj��Y��N������8�C���S�C�$�_|���|[�;�u |�~\�y5"͛&E@.kD��� ���et�qԧ���8�<�*��4��.�9-��O_n�^����꼈�'sz�T�7���(�u@�n���G&C�����GT����4�gw�(|:(�h�E�D�Z��ݨ���'��,U�+b��˵�P7a�}^��Z�Vg3�f�,K�/��>:$��0]_A 봰���3�L���q��?&ߪvb�}�%iDdd��v��v20������%�G���ڧ�{��8�$�VM2�Տ*@�p����$�kFs�cE_pl��z��ʮ�Z/q��M����n�~Lkh�_���7#���6_�L3�3���_�9Û⺖�^g�y\<�1J�ȱ�͚R���ðE��5�3O�#��	�S8�;�ni,f:T���nj���F�տ���mY�n��0�}
�EdPp�H#P?U��X1+	��Nj�o����J��!l1��G�O�^�[w-q떦 �p���C���eB ��k2|����\'�`�b��Oma7?�IS1n?��z��Z;�L	�����W�:��Z!;������N܀���g�`�y'3@&�]�Ε�|�п� [l�X���I!޵ۢ8# �q#���yPD����PR�l��A�]�g ���CCZ��)���V��b�(�ɾQ;�z��Ip�N�J27	����P�� ��ܝ�\���[�C]�>��Đ��~Q�%OѲz#]O"��]#�O��4�Ҭ����8���Xvd��9|�raŜ<@7uT��� ��IQe �"@��^^�xߗ߷���Fl�[d��Ie��k;���}4\��/#��'XR)~ݎ#����� ��K�$���glq�����)s��O�&&&���K��	�G�R����u$}�>�����G�Ć�jg/��b�Y����tjO~4��L��2�S̘������A��c���_9칠W4w���V)N��G*��af��oyj�~���� >��lDo/y��)��dʵR\�=�RNt��S\7��4(Gyf0Q�s��g����n��ٚ�(�i:���v4�qN�0�4��|&6�@L�=ܿ��%r.p䤅@�6v�l\]5�̿�3 ��?�8�չ��;X���^dw�Q�)y�o���=HF�����#|�轸h�[4�fu,��;L��FdB�^��&<�e4(�n�E��T��EJ�3y�����# ���	��w�_3�9�so�DTFXd,�}���ƆNwe�x�%�t�O2�Q���ۮ+?
��M�aDf v;x5ZeE{���=w �xxx ��5g�lp���9�aT� ��M�RQI�Ƈ�r�}����7�u�R��&���C#��)�7A�9�k8� �a㠹޲��m��4I����Su+>a�+3�kʽlɤ����JTt�Nf�0f�-Y��u�bK�a-����UD��
�;��#�Zr�Up�wD��\�D�Y��	S&��,�(U%D����p@2!z���ľ�B�C��x�/]b�֙��j���(#�r;��W�Z��@���1)��<�`�/xGE�߈`O~N�K�Dc�t�h�x�E�J�s��R@���i��n}<�5ģ���"õD�����3�����P�- ��e>�]ls�	�.�+K�5����E~�;�OX����{�%3k4g��!p��Ps�)ǶZk=�����㗤�v$?�"�Q�V�؛rz:y�I���~|��2�W�1�@I����k�"韪P1U<"��>�}߀Td��!��PתN��W�K�F5�1׈*���Pϣ	���EΨ˴�g!�z;J�;�-k��r����dU�v:2U.�ƺ����q	�?D_N�����}A�{ඉɳ�������a��A�A���6����ڟ��7�:^?�lO�T�@�S3Pǚ�|?�^i����.H���z��d�����Tw��;Q�ŖVyt�ȸ�tP��Bz�d��Dl��)b`�iw;�{Q��G�f���UM��nXj]�b�З��dk�I��Y]���X�ks��O����pǖ���7�j�m99� /�ėS��---�� [f�bn;Z%||��Ѝ�x�çCO>U.t`=���<�F�|M��ښi�ҡ�.d���?�҆��r�=�2y�2�+��L:��������Z޺ő"��!�}M��a��\i߱��8n#q�><�����$mjMu��5��]�$�1���z�ćq�~���^Z̿4~7"�����jx/N|�O7ZK��[g�s��=WRx���q�ed�Qo��ۄ[�u���x	ֽ�0PY�ٷ.bT"u+G��`���D&���j�2l|�hT#��s$����l�&��n���T��\����&���K�<������{�������5�nV�17R��A�L�|<��B�y����(Z[\��R��QJB���TRf�6h#>M��mi
v�M2;褋�ܢ��``�A�� 4t�^׻��b�_�6j��q//�-A�M�M��^a�!֪e�3��hh�1���"9J�3��,��7G�R@Gbt,�p�?x�B"�v��Fs��b����G���'����{[�a5OM��1)D���C7KLHh���Sg�T����&�5u'���E���1�����5vI8ť`KK����% \��{#����x��C1�4�����x4z���zc[�J��~dmii�u��ש���*M�[��JѸ��Eqkj�P��Ƀ��x�&nX@2"��p��(._߷�Fjw�� �}�*�3�#�S����5�[��m��ʖ�t/#dc�9u¬7�&��oqKz�X��w�Bۂ��z��� �?�D�ή\ Q��[�9e�U;��η�u�4�T7�aM��9�rU��ر��5g%P�.R�'�|��^���ѡ2��w �^�C�e3*��j�˔�S���V�U����_.�U��sN�zԑ�z�V]�S��sLT4)|Qg<��B�^�l}��y}#ڛ��mGh1��2id���;u2Bϗ.o�Tm�Ib�JJ��ڕ|J�GT�{���z����������_J�#x>08D�����;�~�n�M�$���G�k�I]�S%r��fOn��z��=-��M�s}��娗�]��=Z��#�GmuU%���Q����&]��8��I�@T�;a�i<����K^z#?.�0�S]��/���}��y#���qv���ٝ
V���Vz��då��7@V� 4Fu��)vx/  �՚��������u�%p���V?��u����.���(&��Μ��"������<���ª=Аd�=��[i�j�#/��^��ʅ��;c�@�s���%���d@=��6���S�_��nY/K@/���l�N���s+�*Y*-�l=��H`0��;b_$Ѭ(??hb�Dg&�a��r�mx�PE�7��R�
�7r1>E���LS�q\����.[���5�ky�\��3�����S�X�.�i������V�}j�������'��}S�^��K� �#*d���,���+w��̼E :ⓒ�����k1�����i��'�!��J\�q���k�5�7��:>�\����Fb'v�Vq�p_��y��\c^����閯�K4t���"��V����]F^G>����Ѵ��\�jc�8����������@d�9��V\�~��K�Iۙ;:6���+�v�d��~f�n�P��>*��F�bg��m{��o���q�S�ҳg�9X�ӽ�/\*��g*fϥw<27�G�7���!-���j��M7�^g}*�wP/A�h!
��s-�c�slʕ���1�=`����L_�tp�p�
�_���1k�X����B��&�e��'H�[��y&G T�Ҧ_� �a�ت"A��g2�mX�&o�u�n�����
yq��V�!�x�Y]�'���վ0��a���Q�ҧm�]�	�[��2P��Z"S6t���<��(��@������k����)����͒fyYG�79�� :"���%(e���j��6W�V��A�"[d���?��oj�0�Km�]tlU$ѡ �N���(�bά�;2!l�Ud�l�(���֕ ua�| 5.�� ��s�X��`S*!����������}��H��0=�13��������C���^�0�C��v	�MrLj+��@���w݉���7b&sy�Nt���6I�x�v^DB�A��]��zn���L[�����с5��7��ߊfe8�Zl����g3��O(`�V�)�$(͙7&h�$��j�W��nha`��yO����t����S_�N|N������S��z\���������{���-F�y�b;�� �����P%�4 �[��A>��n1׊�x-�5�N�m��r����Je5ӹ�H�-��.r��Ƀ9�|-UzSe'�����Н�޾=��pP���<"�Xa ���f98|�2�(�`��}¥�ձb��ҍz
(��ru��$�Tu����L��"�Nxnܮ���H���	~o����q���I�u��D�F=�"���-�:�R)h����;zU�w,���l.>C�Wk����wu�@���`�'&V��$�'� �z�4����5;�E�"G7Cͼ	?�9(o8��k�T$�aTE�I���1��7ʫ�6�}4+Zn���9��1��`�;�i^)=�׈���E=~l�Z�@�^�߅4W�:d��G�}+ڬh-��N&� =�v��%s�.��Q��(�#�a�RՁ#>�b�f�s�z�FR���F�	��d��.�)hT�A:�(�bI���W��Ρ��{(**ඬ�/ "���PB���g�U6m�'�&�9pI���r�[�zJmq
�'G��B��̹�F��OrK�W����FB�\�sT�'\�q�-7��4�?��7����c��/�9�=�����h���^+�; �bCC��c{���B�VVW�W��^��V�i�P�5������Q!b��ˠ�ܠ��12x۵'���*ȏw�׭ݤ���Xm��\KO���x���p��B]ʊFG)8[�њ��WA�w｢'�!_�,ڥ�^�V|�v(���ϯ n����-��%�/tV�s�`:E�'��Nm��W^�b��ҥ�����h5����x��|.�j�{ls�V���!S���'Ԥ�ٳ���]����'W����\�.ߗ��4��kZ?C�<�}X���MT�F<k��Yt``��8P �MLL8��S�*j��4���SC�����˕kz#���p���E �0��FT���l�����+�Ic���?�*���a�E;=8J����gAH�҃���݊ļ�(�b��ɷ��n8����P��T��B���<<�b�~(%�%��3�^R��B���3|h������X*��o�׊ �pj%%}��n����0�'��{�k��=ș��D���Bod���Q��Z��L5W|��������P�j�6�CV��'7xF0�cG&�23f�<5�c\w'�@n�3-ND����s���8��F�X��!g��Q�ŵX5M��R|8�S&#k!_II�]����0#���#b�����Ĝ���q��cH�f_I�:2agP��#[��^�9�=2n>W��j�,L�D���稰���:��VC��+Z;�O�%(����ï���{� n}�N���·Cte}�F0Ӂɵ���E�=k@hٙ��������@�`�C����I~�%bZ	�De5�ӳp��j;1�#ur`��)E ���|fR�B�¢����"D7ٛv��G�����f
� ����e�շě�wҬʥ3�h���|�����^ʥ�8�A�Ѧ��K#��.�g��������Z��w�{�����:�l~3Dc���Ԫ�����?ٳRϗ|�0>�^�f�3�^%,�6{Eo%l���5�3������O�b�Xk;;�S=��s��s���zj�Z,��z�v�"r���G�����n�wq
�C<W�B���c��u��H%3i6bHmr-�3�m�j	X�?��4}kB�M��Հ����6�\c���G(�3�A�	����`ُ�0}B��ڌ�ho�^�z@�W�׵җhO��c��g0���>t�3����=�o��ɹ�fn�iTL��ߝ�N���Jn���@ �#p���<�h���Jm'�oǮ4:�X|S���C������iy�Ў�]]mP���!OMF�t��?s����+.=���uB%����:���, 1BY����q�c*=m�M����,G�j�[d���z>-�-��]�\]�3<���񛝀���rmWE_�Z?5Po���%ʷ9�j|6��|��"��ѽ]�z�^P�/����q�x�2kTB}��!��	�H�h�=�b<�Gc'�'2�z�~0�;�0����[���Mm+e�{�u�f�U.=��+;⻟�%2�	8��+++�{~v�2@�u��QO9eU�4e���-�==�6� bv���0�����V�٣2���1`���3i��#H�!���4�Z���6�(����)�֤߽�8���8A2~��~�j�o$<����81FJ:���^"���[kT�����,�����E$hr��A����% 5nL�*$���L�,!G�V��XD:��F썍��6��IW8�Ӣ�H�AB�]�- ��&�Rg��6�0��z�s�M�z����w*.�sk7WD*��t��Qd� }����ȗ��_��H��G�+���׈��@���0��޳�<������j.6]��M_gg��.�����|�ӵ~{��/�ܖ�"*ʌ�V��E!��m���-�7�O��w�&�4܆U�p�0Z��� <�ke�>�i	�,�[��gkF�qRd��]��چw����]�_
lq��90����J�=0^�����^@l�:B���_���a�ɞY�n�Z�"�Z��3��Cm��/����C��
[3��ː���MO��M{{U�O��|3}�t�n �8c�՛�eUo0eB�t��d�NK��A��]�֤�&�1g�x�>��Z@��"�`�hgUT�����Dúz���p`xi@["$(��6i�+)q-��3���;w� Ln���+/�Y��I���{��r��H��5��C<=�Yf&��Z�ͬ�%��{4Wp/��6ƽ�������$Da��a��IBc����5�h������^/O:%R����I`�j���֜��zz�5=9����[2��l��=̔�c���l����d�}�#.�x[`���>P�Ga�l_�#S ����9�
��G�{�*��`E���x�^լgO �	��������nb�Զ��Fм
�f���dԫ�	��Y��"��G�Ɋz���$�Dtj�w�uw�k%�� 3:d���Vy6]�f$�/���o�J$%� )S9��}1((��i�$��߯�t��=�2�XGG^ri;M߬O����[n��a�LTe||�`��zQ���(�S@)� �4��v��Z�u�����'�ydJ���4I��I���1�>{(T���H����q��x��Un_���Mne	�M�k@A��8E�/I�~x�C}>{�,�m��"�X���B<�29(�>@N~~<2y�o��^{e�(||`o_���K�ug?�oT����oHO�	� ��D���iNe�c�`��vuբN�����z��nKG��#M�Բ7"�|�.���t��]g��3؞5�
E��|!#	���ۼS����_s�@r/V&���ܰM����p�u���#+7�՞�(X�`[�㜉�	@�f��!v���q䌺������ވs�=�l�<��5}��Z���'^��6l@�ӏ�ٰk�HX��TT+�x&��Qw����RS���2w�b?�d*�.Հ�Cl��-Y2�{36(��Mzz�?5ï�u$O�[o#� ��� 7Y$z�:6��5P��i��5J
�>���%�
�9I�y�bk �}RNh�G��l4��:��R��e��C/���Pq_p�����i?�����Yu�
T)r9�zl���� נ��������biY�#�UX��R붇���A���D���3򦍒���@���I��X���-+Fߋ2m�/I�U�=��	� ����	���?�r"Nkg�0�Y���l�qR�<�{�%�&oU�f72���Δj�*��* �^8�+����}'e��R<ڮH�ۻ�c��Ѕ��l�ł���o�īh�Ǖ�h���Aq��_�4���r���X�;G�\�v�X+�n�}�$��84
vY��1&X{�t�@�R�!�����~QvK��-����h
�=���C���@K��FPJ�<���BZ׮��_��O��Yԓ�k��c����n֌:4=��hd�O���V<$�äTop{�G���]њ���rp	�������I1���VO���(��bˇ����9�N>�#�k,�w3�6�>&^��p��,�3X��@�;-.m�A��DȚ�$�V��.��PŲkW\��W~�A�庠r�*Q�u��f��Ml�ºE���IV�ʈ�̑Vj���0�3���!��l;S'�ZMS�R���j�OfhV'#���<��}�\�l��m���oC�l�����r�D����+��-%���u�o�~�ݨ���~�Km��ş���=+���>�S�7�b��7��������Nt�[�<�ǵ'�+��/<����P����A�2�X���ȹ����V���?��6��,2�U���r@{"�v��/f����#ã�Y vfZ0�#ER��f��`�qk�<���Kq�� �
^��mju�������׿W�VYw�\�e���Q"�o��E���N��4\�Wt���9e>��&�_�I�N��m��V�wz��7ʓ�w<�g��;q����,�IE84�=ux�I=�����Q���8��|Fl��@�Mg5RH(`�Qe|ʶ����1}�'������C�� sKq���)Ɛ�м9���Hبk�ޭ+���2��;��!�@�m���X�)7�X+��#ރ�T+��-���an}��z:�������ig4���VQC/૩
��+��/��Rq`�O�,k
��6��[�OYk�i�d�e#���ꞻ�͒���&�Z�"p-���!̫�l���&��ZM'� $d$���D�N����w�".8q�Q���
��R2�G�!<#�E�A'"+��ǐ��N�٨��%��L�L��f3A�_��NO��?50�/ӑʢ�lm;��LT��]�̷�5�v�Jس�N��Rc,>*B�=��|ʀ�R�/�-,��j�uZnZ_/�J��`_8l󏊻k�Cu�O��UOJ
��H��j��]�����e>k?
Kih��"Ǵ8���ɅV5�i����o��{��n�>��O*��HР R��BS0�������!���߳ ��)������c���C��-���}�鞵�ؐV
�1H?W�䁶L���i��g����0!���!#ǲ6]dJ���z�n�������٣�$O�Alc{��P���f��vG�����uš����d#�P�
5m�w��h���n�U]���a���k��~�3���Z�N�_���=bE�z����x�WO�8/�� ��l]t�@[ ���T��3Kٯ��.S��<e�������JD�x�������48�uO;��!�?K�{��wn~����PMٓ��*�\��Xx�vR$�kYw��x�J�w�&{w�Dw�(+O�A����>�m��;��q1�j�(��{��B�����(���u�b��Fkc��<�Vhj�P%�z�[/���A���ԋ��!�cLw?׉S,0�6o[8�����n͒<�� �~�.*�?`�q	 +(!�����������>ņ"sg�?e��N-�/��<��}�[^��F�P�3��Tz�T����٠���7"�w�N���ӻvǵ'�i#�GJ�H	���_̳����V;���R��^#��4�0��Y�H�b�vv9GohU�?�7Ɛ;��Ɗ�F��N5��ߨ�sP�/j� �ķa����N4W*��X8t�ޱ�x>�I���m-��	Q�J�={F��i? \��Hrb8p���e���P���`K�� k�[� � o ��[� �g��@aG�^�=OΗ6�&�9V�̼(��/Xb��_�D�:���ݳ��B�hu��{��~>ɷ��2�}e*l�W. h<��/@��4�Q���ރ�耂t�j*�n�L+����n�>y�\�W�j���Pzd�cnsC|�>���:���-���p��'҆`��鷏���_�C;Ya����O,���^ �Wff��Y\��D�PSYlHn��V�C"��A���ډg��:-���:���9�k�ٞ��oj*�k9�	D`K��N=����+�����x��x�:������4$.�iL��_��/&Y�U����S�����F�+������t��6����m)����1��>;�,0�UXRRK"���Y�3y��Φ*��È'�q?ל}�%a���,�}�=]-���YV��D�q�)/� �<
�|:&z ++�Vo��<ǣ�-�p~�����捍O����5�W��i��C͟�X��~��赔T�i�N���s��ϟ��b���䖿'b���'p�@A�.;���:���m,@AS6_�/XY^V�8������ox��o����*+G����Y�C����Fs4��߫�O���{|� ��"�zN8j�#�{�P�����j�}�F����	

�ON��F���,������e��͠<c�a�;+�!��_�� ��௷��L�������\��*+�Am)���{�/�'���If檪�����<�H�spp���w07����5���J4�k��F�YY�v��������������:��NVCqaaH�إ9j���(���Ç��]w0hOmy�����ݯ}����H�,//�.�GB|���e��!|���sT��Q 	�	�����L���3���N����   ����h�hKuh�!~@-�"��\ o	�엿�P�;6V��f@EG�FA(�m��es���('�XCK+$��,p�\�AAA�#kDw���^P��X�&gUK$�SQ\A�����ܯÅ���hmƲ�0��?��r�`[W�8gp��37���C7跞)p�����U�����>���γ\{�H޸[Q��v'��oj����o=��wS��&�������=�n-ߔr���"K�~�bٟO�L����;�s�����W+�@X<�i#��9�P?1�N�cP8�*���6��n�� ��/�q[�l�b�_�]�����<�����54���~����,nթV��X�s[Z�V�+aj��T�<W�S��hv�%���Y.�'P��������L{�m��8ׄ��yDm�/9�\��R6a�E­ixh"��5}k�̰sWcB����f���ס	[�t�Ԥ�%7$�4���4E~���9\�"-L�K�h5u �j��9`�F7&��3|���0��v�ױ��Nv��cw-�����q�I��~Rҕ��I�Q8��v{��_^	��x�BR��{��L�$����8+�����0�u��e%��`�Rp����zn�n�@E��eG)1m�������i\�#��(��6��@q�ݥ��;��R�O�Ȩ�l4E	�ye�]4��1V��Ox��E���m��2y�(	S��FS�� ��-v���,�z�ܠ�H��_$��)� p˅�o�����w����	������b��)"	��E��F).!b�y�]��O�u�=�#>G�);�S��5��:�I��c7d��m���_��η4&{h0���w#B��:l����K��<<<��� }�4srr�z\
�ܘ�:8Jp�LBId-l߭�o��>4��\?��K�$y�����8���P����j��t2~�NG>�Q�"��<�����Ԫ����G>�g ����LjFݳ�f�xC
g:Q���1{@�)Y� ��6��,����Ҭ�x	�h�C?lg�7j
�TNE��8M�9���ic>Z%iT�D}O��J	�9��ތ�]����t%�۷^��K@kxt%�>�
^*���2:
��� �PmD
����|^��b'���se�eR���'�Q������0��Y7��]<He�ڶ��%K�L�T��۟9��ok?	.(ѯ��_x_9���h�a~��-/�V�mޱf`���9���Ƥ�xp��@#-���k���4�Ż�ѿSU��!���R�נQ&լ��\�Y���[���b���{���������+/K˧�ۋ�@� ~�{���3� U.ܭ7�qY��e�M��}���#�����Pb���/��պ��5�4=3<�1�^��E�ZyTKD��Y��k�~E���8Vk�\�dg������
�;GR�"�:���`Q�{��*�v+�w�L�N�����DWJ�4iۭ��j�J�)�1��0�j᧥����~z+��N���KD&rЃs/������R�j1�N�{s��K)>8�Z�g�������q�J'�W!�KB����/��UXN>V<����ɸq��P;�:%I9%�i�˪̓0�����r�G�F���7{5Ggt��n��jH�|{�}O������ ��g7k���4TUo&��^p���U���w�����D������3f�S�)���/�������k�B�;����f�<�=����0�y�3���w*�{�vZ%��������>�\��V?+{��5��򇲘��jhzl-�������2�d{�s����y�uޣ��|���'��q���,Ͱ�f��j-�Ct+�RˢU�����a�Oz�$<���R�ec�9x��0偬c S��e��{_�R�?Yb����I��3�I<=Z�n`Ps*����] #���(��u>��E��zS�{��k�����NSLq�텛�_=��zs����w{��-!!q�8����dk��'��|ƶ�f�e]�b+���)�H���:���է�S=""wF�����[߶��?T��j�4�Y��u%f�o�K�^������<��t��q��[���!S�E�J�\�Ͽ�����/�����n���#�R�ae��fV�BEK+H��ԝ����������0;���['���^%B�ʌ�G���>�j�ϊȬL�ACW����n�wE]��t�nѲq�y���/ɕ�"���wŗkh��EЉ|N	�egUp����@�>�ק�>�����w�Q�8��.wETݵ�]-p(3ߎ�t�?�x����%1�ؽ��;,Ȧ�x��f���u���}+���t�9���o�]�JW����ۙY���tt.(��JQ	a"��Gl�%�a��Y�������+ (�Ɗ��T�]��R�C?�9���|�]�Ue���nz����k�Z�9�S"8`�-�8�%�Y�z�����y�B|f{�M����[�M�{Y�y��9��W�e����h�sAfJ��U�Ϻj���D2�}�޽�A&h_�	
���޽{���VQ'��ic�F���_f�э����O��e;��^��#�Qq�9�)*�V�����C��,�����c3^P�/�
׸跻��dO�Д�u���/ɤ�ۚc�=�6U���5ut����U�H̕D!�ּ5b3ۥf��4i���y��k�ќǜK4�7�`�E����P��mP��fpT%�������	qu#[d^������ <�� ���c���!�xz�������:}���~�ue�y�B�c�h�o��
�g�������r:x���ZvN�7�s�E�()�
���b�����s	������[a�"$O�kT,y���{d1W)�)�Ho�d5ɉ�5���8�ZtZ��mf��[|�w�Ia`�"��;ˮ��'R�m����'�7'������6/�����-�e>���O������P�- 
�jrʿ��^K*:A[cQJʼ��D��2.�JU6�M]QJ5eQ�#-Q�e�Dԉ�e�.o5���;r5�!������W�o.���5\���7���y��$��^dq����ʿ/����*$�ɕ4��ҷ`uu�)��m� ��'���+@���.�+d���DO �	]Ee�*�Yi��G�������i!��r��ȝ]O�Ŝ�����Uei�a�a_��D���d��4d�^a?A�#h�b�$$�]XR"}�i��r��ůA�2S�[oO�������Cg��qF�b��
{��m��:2Sζ�ʻW�V|7���{T���ߺ9S]�#L!�9��-^�*S{�>��j�#����0B���Ĵ�=RW�z�����O������dɾ�������O���,'�f`�g��m�U����{i�����\�x����EB�)���9�Ⱥڋ0�w֯���3�Ĳ\�c�f]f���	�OGy�<���Gh�<R�|��_�ȋ��,���47�ĳ D�@�m�{�}����-�C��ؔeZ��a�'6���ڒ����|Y�x��
Ӭ�| g�"s��j�8�������8O�L��ޕ�������i���iH��8�o��E:��W�#�Yd��&��=ʵ�{�15�I������������ª�5��SM����ݻL�-E�� -�{(y5s��%��zC��y��3����b�Ɠ�V�ד/�k���M�Dڴ�i�ǚ!u�WDu��u	�察
��i�t�����ۻJ��(.��=��
��o�H�(R!7KlR��4�p��t{�ɞ���[ݍ�<�Pվ_��em�f����6"�XD~>��k�9@��prp<24d<"|%�BIy�K��
g�I��~B��`��\���~�eE�U<Պ6����3ۯ�c�'t,V�o˒�|��B�~�v/f@��^�1t�rD�����\ĸIx3Q�����e��?~J�'è.ob�r���kʗ�\��Mk�x�b�@��}�G?L���11ީ�z.��MK��S�`���7��k��K?Wz,-�lnA\;Q�:��O�ͺ������IaJ�;!B��׏~=�m��9�r�p!%(��Af�G�Ї�&�W�'���K>�+ڟ�zPJ&��x��溛�#�Ȳh[E�[]��[�7�i�TxIik���[Vk��$�e�A���Q����̣�o�-]�=蚎f�/�W��~��={4�y0by��(5�ğ{?����}�I(��}�_KfY��0����5�
B^ ��c~>IJ���CH����NM���MY7�yۉx�cj��̄A}�Q�_������!�xJk;�u���%I�R���lH#���D�Y�K]8��f��C�|�9��W��e�v�6����9`L�X��L��h������b �]�	R}��o�6z����U��R���Ϻ���yz�"pv	�H�ߠ�485�ٯ��敤��8xxd��%�^�
��#'�[a/��Ǵj&}y�lS;��L.b��0���sJ�l��FImMO���vI�>0�:G _��-%}�G����'mY)G�9.��;��hM�Ic%��&
T�P��m<5��V�D��d�M�+�
��~"�c����{|�w��,-�Î��[]o)Z����)ۇ�$�<��C{���y�,n�� �R���-��*P��/��ԥl�}���^��տ뤪w�����y�m���W� ��v���j�V�����{!�jg��p�2EE�o%zu�2�
�ߖ��й�"�5���3���ƜI��Y��
j��ݷ�|�N�o�U� ��1�p_;] �������L3��S�Y�)){�m�U�B���1���ju���V�)���?;8���~Z�٠���\@ ��d�����܏��.`�ZV��x���\��_:��k�����jh
�����CoH�Ժ����uh(Y'�pc�顡L/!J�)���5v�����cY"�[�4IS��%�^)��6��3PL��ͼ+ۢ��xP��?��׵���z�1�C0wA��lf":����Đ`��9�QW����S�R��e��9��ش�"�L]P��4�-u��\w�#� L�2��T��$�k}��X���i�Q��9�x�����/�g�-/��wtv>�b�I�#�FcD��B���דfwf��vQa�NS���"������c�=��-�f�
��bX��� 5XP3�	S������w�Λt1U��M6{��NtHH���d�z��8(N]����/p��Z-�.?̇\kT��2,s%#0�i���z���l����N��u�+W(]�ZV羸U'���1S�w��R����xa��]�ОX9b�(L	xz�3-�Z�:���=��u��3v�E�P�^i�|t˥g��>��K_�8>����#����=]|���\��36#������9�����;N�O��X'��,���c��&Ů�	#_�(��;~�A���p�Ж5}���~��1	t<����2!���V��%X%Z�bm�GlIn���b�����ȳ�?N�X�-��k��Sqñ�ۤ����*��:٤�b�Μ%��g�!���B��9o��Q��lR�I����v&����#�0�������΢ϋT��(
����]�'���W�c��� #s3���gq�7�uq�(����wUM�=��'�E��`)���������긨���A�CJ�F%��TJ��;��2�P:F��C���;������?8�}�^뉵�>���\r�z9�g���f���0������,�KU1M�X{^|�k\������~�AL;dTHgb�����/�-1�N+�~�D���R�F��xK�};��ײ�ʰ-3$<��NL�rz~~U4��_3�Kwމ��}~RC���7�w� ��?����k|,�E���	TR��pf��r �K�}EF��wQ-*���F)��lug��K�܍�Yat�
�8�LL��]>�� ���G,�x���߂�Z@�<�4�9��W���]����8�Q��0��I�����U�h�z�؉7`����\=N����M�5Ȳ�]rh��d���PYT]8q qp�:u"���>��N���}3b�|�S����u'giG�&I��Z��}ȵ\��b������C�:���r�����6s�؁'Y�bA�i �6	�Z��W��<���fo.;L89�ޗg�?�yS�b"O�0����'^[WWn�E���j�EB�F�����	~rjhxE �s*rb��2�$k|.��{����b@ԙ�r���ҧ}��`�i��xG�&��#_Q�x������|�B<��Lg՟�Z�����	��8����(����M�)��!�Q��ch�z��:7M�ýp3j<���x��T�����W���+7���j"��f�W��m�W�\7��m7t�����w��Q�k�$�v�7��xY�HA�tW�˨Ev��HCu�[!���#���!��~�+��eE���W�=�j���Q՘+<�9v��9�� $?�N�v)����$���A�����ŷ�&�jq���N�s�^���t�Ղ�z`u�Rp��?�=��S��qU!��{Sj��e�V�k�A�j����#{`��_7�r�هA��ά�l�x&R�7 Х��U���H�pOC����X��t�E��ן_�����F�Z���/���yыɟ�3E�=�����g��������D���rȍ�N�p�}+�3�@�qNif�Ә��k����*��v�"�#�d�!À�+k��@9%��¢����G��� �nǎ��K�%]OҒhܰ]v�ClLI��9�UǪNPd*�!�	f`xo����)��j�ow)�}�0Z������������`�G�DZ_|&���69�`ܖ�c���oԏ����׮� x�ʤ`�����@A��ϱ54�����R��%G#��­�S�FE�A�����'J���b-�a8ڸ����Y@Ff�)ī�{4�.y��|��"iŹR�c��Jm覈�N���ؒ��s W����I9NH�e���=��SW�r`s��?�$�'�Irer.�,��_����IiiQ���ii�i?�p�l�������X���W��!X%o��D��["e2�	e*$��K���w��G��I��e�t��z	BV� -�j[��#*�$��uZ_����0���ݕ�gë5R8�(�UL��j�(�?�I�9�Su?uf_�@6(LT}�����E��op��b�e`���2��q�E�ޱE<@M�5����� �k�|?@��8���<J��ȁI"���D6g`����\&}�W^1���X�&�Wy?��j��I�z��H�����9�T|�y�y<�wVd����Mp�dT��=�!f߬똨
j׈����]������[n�G9�ͣJm�lr@��A)a0�e�Nu��H@���LV����/F)N
�
����բ�8��׾:$��!E,�����Jז�ƺIݯH�����閄�I}�⦷ �t%]���n�dj�%�&���=!�n^9Zʉ���P&��g}�|-K�[�@��+��I�=?l�V�1(g����c`/1�L��󽘰�w�"��WM��1���[DkJ%�$��g
a/P�6�do����b�u�>5�a��*����~T��a�ogs�y�ʖӤ\�@JN�t㐂v�+��ʤ�h���A`�[4�9�M���đY��]�!)����P֠��aϱ�T�4��G��U "���~z�_�`j��@m=����]z��c��;��ǂ�n������)���hh�72��Ѕ< Eы�	�4�{	i��x��$��+����V��*r��K߾�-�'#9�Ÿ�?	������H4����DQ�5���mf5�~�tݶ'n�XiF��N�6�����lR�)I[Z��]���������!*���~W@i�@ �]Pڇ)�'I-�1:Óh��WEK�.i�WZI�>#?�!�"7#x�
l5U?�J�i빬j��2X�{ȟ	���i�N��>���T�a�@
��֓��1��C�T�ꈦ��nZ�y��p�Wt�����C�:�YYh��x���X��$h�d&{�Nqw
�RtZn�|��Mv�UvC�n�"��H�'y��������@S�uJ&�N�[-t_�x"���"S�.U(�݂?-���W)�mn�����������k��s��N������44�`��Gb�L
(M���I�u�'����7�����cn��fD�zVM�"1q�[d��9*�o�dA}T����B������p�nu
�d�*λ�ºո�M��1X�����!��A?���W�kb�&�``Jɝ�M�ZO2Y��'����[j��]���>]�m?Lz.��&N�*j����Un?+�]�Y�BD��?���O��X�u����2�ֵ3ړ����}��ʔ<�����`P��q�q?M���)"�G>���9�}��$L����(��Rz������7?Yp��cp��C��`�J�`'*K��&|���|9�Wd���ٽ��{���]�C܊�Q(�e�ζ'�M~0������:ܐ7��IL^^�\S�����8�Z�Q��F}����i)�p��qkLfe{�g!��sf�tA�D#�g�z<��#���b�u�6�4��%%����� '�c�ꍠa�}�@{��^�D1G,��H0��a(	�Ltr!�s�z��*��"$�c8��I�'&<�H���iC�iC�������f��g��j��\l-��YiC_l�=P�FSt�P��f���	��f�!�\o�����ˑ�p���B�w����bl&��VT���\6�\�����_3O6(ZM���K~��+-�P�C��g�|itK���^��z���Mw0ڼ4��O]�O����Ǔ��� |�Њ��E�I+���9�����eZ�W�­���V��琏�T3tќP2�Z�;o?�����5�D|��̀��#��Z�\�pp�0�"`�H@����RP�������W�����e �jz�$��!Dt��X��e������������>��:n. =Yax��� �����n~�P7=,����p̄oU����� �?�#v�?����x�S�K��ǌ�O���{�P���W��|哺&VO��:{"�s5i_��^8����s}�H)i�p��1��Ƅ���n�1��^��������ff�O��%�� Ҙ_��)���V���Mzv.�Yh��,���}j	
�Nͼ$��)��^�qM�Ɯq��<��-���*>HbV
�^A���잻�D�b)�I�8�! i�X������s�,��h��}ʸ:��`�b��W�n��>`�λ�x�8F}0ܫ��Gy[Y��Fs9y�-6�d��@��t7I"lDB�0k�
���E�Y��;[�&�3�m���/�0������=LǱ󢹚S
O��C�'UE<َe>��F���UVr� !��t��wT�l�-�X�1��sd��Ao�MG�X!��r;��le�&�3]����-��&:9c�jD���Yfi�U��B�r�%����o��K���^Hym/࿖��� 5yZ����L<�Mt�h:f�xh�U����>�ӣ��]���Gz2����8���;T:�j>����Z��ޫ���

n8�gffTc�g�M r�9`j�/5�*�;g��,�^������%�n��#ב���Yg�4�f�]���\@��}������w����F��9d��ĉ
q�����B��ɤ6/2O�@:�U?���I�4in}��0P^�S�����/��/��G��Y��+��~��ZΥN�A�X�Q�˦��]*@�s�o-��וNYqd�sAE~Rh6��i͚�HO6z=K��p�d����v�(�US���2qܷ����Mw�a��O��g��j �/p�4H�7��d�Q���r�l��Zo�_�'��v3� ��m�@�4x�"b����j��<6qr"r��~�U��PGZ8[�N��4a��P �� �Y�#�� �n�֮��Zg�����|>�~��q�7z2�d(��EĆ�+c�{�ړ5=�'�Q�9�3I�w����-Tb�=!�x��ĸ����s��w��-hmܤԇO�~a�Ff�&6-�D�(��"�t�m�wc/�2jj���^6���y�G�dq�po�+
 j~�q��T6F�=�(āÞ�!�g8�O6����I��c��_�0�L�Lz�X�˲J�[�e���2\M���aք����Өyt6�6�Ǥ�[i��c8�j�(0��x�@~6�M�2�}Q����hJ�ƺA�xĊU����@l�θ1���g_sG�UMaPq��s��v�S��G� +�]�/o�6w-��/�l�|߲?CJ�4�}w*����n�C=Oy����eZ]_0呐�;c�Vz!d	B��Xfn���3RyY� ؗ��a�/��{֜�fu�%�F,���Ђl�I���;3��	��~��������М$0���W�Y@�sB���rcst)}X���W0�����s,ʯ�䤄��# 8�
�����췳�J^�7�2X���!V��Y�mͶ�v���X;: Y�����a�떵P>����<{{��e:"ޯ�'~�
�	I��K����zڳ+T[<]y��r�G�5���D^:F�t�40	�0k���'WK.���)��;L_�J��=K`Qz �J��ڃ��
����xA5��r�Skv1�����bԇ?�v��IW̄�*eq�����tw�b}Y��S�o �_���]?��}g���@H����{��A`B�	�}�S���L�K���
�"�����{�����R=Yr����ԡWoP)�Q����/�Z��.�ݲx���HB�%
�@��؍%E��ӄͷ�.Jc �����X�|�vy���w�r�a��c8����y�&~/��l�7u'�S]*�%_���MrK���p�r�zLe&z�Dׯ'���Y��=.))���j錦6��A�� $	8��;�!`����=��v�`}j��J�|��q_Dla�r����s��P�Px�ڸ��#�s�e�:�{%#�	y
�mnd��GYD�Dhm_{ٞ�9���<0k�J��M�)j�M��`�\�����e��HA}�'
��ĺ�2xhN4W=���C�H��@�����Ty?,o=-�h�����+�vY�����-�8���ҊT
���Y��G�����Dj�/����?��őI\�g����?���&���ؗ���X�/�vP��u2����*�;&�xx#�� ��c�S,i�R���-�o^�n[CY% U�S����WYm�=o5��
���-�Ơ�B���3<ե��ԝr�Hf���������*n��M�1nv�*c�K_ˌ`�~jީ�#Eޡ�4�ƽy�����t�C̥�c���5�L��z�C�;l�7v)�n��&�վ�_�w� ��(O�0P��P�h@�0B�o#��*9-8��1�F��
��l�ʘ�5m��un��Fϯ� �,��K� ~l�C��[�?[VxL��n��q/,����x���~���!��4����aW�:�Ô�v�����X�� `a���-*��Uo�? 4H��Tr~m�h��v&>ea�b�-��3�fF�F����Z�XV�2O�F�Q����,<> L��	�o@�&�'/��6��S��a��Ao�>��6O���oH��І�W��o:β�x:>��Q�>�
d�4�d�!$6'����䏌�G+��K�h�?\}Ǘ�i���PU�H.۵�����>;/z,�|�	�V#
��=��M��a(B�q?u��((��Z>ʫ����/�3?%��,+{�T��9�1�q�.@��{aa�����@�2�"��uCY_Ai@j�������=��z�!<��4l#/T$��}�^�k�ͣ:W.ÇJjo?G��b�=Z�>���/=nWv>(�p�e��R"�#��O��\i�E��*d���5M�q~��0�����o��̪}O����MTQ�w�t�L2ϛ���Ƴ�]DٲR��H*u�U���D�Kl��P'���+���鎔L�N2 ��Q�_���I��%~�=��L3���--4��9���GAA0�?O ����t5�k;��G�qTK��^�k����b>Sܥ� ���2s�e_��Gw[qrr��oO9��I|6���P#��B��!���{cc��h��"��o�^L�!�1�x�6��P�r-�nʭ��/�^Rs��`0��.=8@빴((�~\��IVE�\�ͳ�/���eƸ�^<�n*3��ڏ/
޹64H���d#�"Sw���w��p}`=�^v4c��/lohWRP2E��W`�T^�c��D�?�`�.���]�=�g��48f�����S༂td*�|;�!�s�ykp���M���=�[��"F)�l����"��8�@��*�i�u67��5�t�.�}���8$DK���#kv1�	b����GKB��~�mg���&��A��csF~*	@,cOj���L �?��Tʡa�+Vz(h���o����r���Aj�����>��M����R�_��^E͑[Jy!N	*;Jd���	�`+� ������3�_�w��ޑ��eH���hc�� 	���Gi9�&b���WN/�j}��Z�����SJJd��u��#��ih�/
�5���o�\s�)��]��7O�Qx�l�>��{�>y��hn�@��؂��?����w!N�~+��F	0��d��<Q~x��n/�  �Il��
'�6,t#���O��HQiF��yA���p����T��SC�����P1�M3��cG���V2�q����/�w�FffzQ�:��ӭ1�x���[IJL���H��A�ݠ�̴�Pt��x)�x�9���E;�_�����#ޑ�^�; �$�!� ]�f�1����{nM�♊�#pQ�P�Z�3�o�Ҕɘu'�a��[�X�B�qǟ���v�~��B�T#��E=E�i�:��� �/`�|_�#���6�>�����(1_c�F 6���2c��vؼ`nnO�p��&��r��\X!`�޾���C�hϠ� �\���l�^�GIt�|.66p�;�x+鳕�:V��ĕj�	�b���9o����ﰠ��޸
0/�k���U�0Y%粦m��dT��Q���N>��;�J�ME�+�}���ո�S�/ՂJI�h{�������t�����J�x��G؆On�����ҟ��\Y�}���/��NvZY���cTv!GrJ���|tY�5.E$F|��)q��{���o�p$�C��	��Ce��̻W�;t)���D��1��ґ:>߄W̖����٭��I^��U���!�_����D�d��.�]U��Za�5� ���H�l4Тk� ��/���4N�tA����U^G�h���D�_�T��,��(��;�3��O�1�"Re��H�nn�����a��:�TY������=�_��z0��YT~C��<�8~OFN�w?�s�� ��}.�b_��]�hǃ����5��ZD<��!�l���WUx+�t�Hp��D�̌[�#<��L�5�����>X��WJ.d<�[� ?���TÆ4Ṃ3f��^؅}�B��F�t�[o�ܾ��:aQ�)>Ⱦ̜�Nyſ/4�A��q4g��,f�P�ł�# IL˿�.�<33��w�hKۅ�/�(HJ�l���$��͇�8o/:���S4�`'*}�sWlY�!!�����o*�z΄IO
��-L�U���kBQ���Rۦ�� %U\��U�������J����q�_�����A��0��"���tdc_�=	5l�	<��Pa�h���Ât�b8��>�/�2z���9XM����e����Q���v��M���L.d�@=����4`�⮮}iG/E�5����-S�/�� ��h��W�v���H�\ �)a_�9�7<W4
83���;:�]���P޿A� f��ޙ���`N�瀩�lo� �����[�lPb��$���-�����!qbbZ$�ߔ �{�v�,I��#& ��#e��d .��]m���FȄ����z������/1�G
@d4��3 �(�D5}wq�SE����PJ`DG}� ܼAl�`G��/����!Nv��pynv~��ذ�}���gn�Sl2?-oO�YAgO��PP��c�z1��Y���N��A�~˯C_���&�?=1rh?��"�H����]���v�FOM�L�\���_�~5o��E��=����̢�!��My4 P��ֱ�$��3݈�B��"��O6�<jڧ;0ѣLv���9�qC����+ki��I,U�~�ϡ�6U�ܗ5����Exݵ���V��]?U0J@5��d��;J=��:���k/��M�<`?*Cd�,�k�$0z>�b�D��]*k⽃�" d8)�!���!�C5X��<'V�����n�,��f�BQ���0�~�����H���=uAzJвnXzŴ|�c��p*�)>�_��.׾�Che�r�v���Tl�kx�<� ��f�s/�Ũ�3C�ݾ��ւE�+gt8{A�R�h�*It(i���$�1}��xm@ʇ����V,����>�.@eL"O\���F�s�8!>��ϜzDѲG�Ee �T�S�������^���wo�d���=?DF�})i=����J�y��N{�������u�_������V؝#�iC*���B���Kvq������.lǨ/x�_7@Vg�j��tP��s��p�/_����M��О�܍G�K���1��ė
��5�� �J�'Z���?ܽ�4�׽G�lx���A%)ˏ��U��H�9���W�G�.rh���9��>�9�� 8�ǡ���b�Ε�D���c[
Hvܛ�.��%�U�����{<^:o0�����y1�����W��	�>����ͼ���6�-l��5����;6��6�U�D@7r�X4�ڪi��M�
CV ����?s�ܖZ�qFܻ���d���`#�(��Ξ^Y �~�#�@�q�#��X*R�AǞ1�D�^Ķα�eP���@�cf&�Q�D���.V��`�;�E������'~�b��ܗm�����'�o�^��I��yx�*���Ȕ���=�ѳ�}����Q'����j۳gP&��\�,?TC���V�RL���+@�d���-�\�_u��T���*S�w�6�it���Y�~d�^�?g�5����}��o�ɼ�p^�rm������;P�f| ��0���i�D���qr�m|���?�1�;	ĻRMÙ��3���XU�s���J�������Q�ß���ˡΨ�1��H�����1�5��a�jN��F)���7�,5GJD�k�d����
  �a�t��V��.��CS�zrb��X�~d[�3
 .��<T�(

#J�jL���ۨ�ԕ�04��G��w� سl�qzIS�w�٠�r�S���	��M�
}������R�{3�hf��[:���������h�^��������0B��̒7]�}Z�bM-�K���l�9�#��G�O�%�Mm��]�_$n��1��.���:f����:kj>���{U��\�vmg�I�U�ؑZ���ğ�<�6 ��k���DOk�#(�;F�] 	�:����Z�9kK(��c3-��|@��5=��i�Wm]� p�V:�?�?�����f�G~>6�E��]e6����B\�)���b��\�Q��k���t��X�k��'�	��� n��&�&~2u(O�+9���&�qQ�����g�kJ~|�s
��2�VLf�ש�֒�ƥ�����Y�?S��B��G���F-#��X;��~7O�T�7�d)�����[���o��C���
!ɱXv�љ�!I�J�a�񵄀�L�Э�;&�	�"Jw�g\���b������I�ܴ���vX��Kg�&U�̇,�{Q�lN�Ԍ�X��{�=�kx8O4�d�/$%Z}���4�a+���]���|@:D��<� e������z���:�2�=!��S�co��|&SO�+�
����XUmrhSu�����.A�6FDhA�A���"e1�OgwZ_"
�3p�\d��|�_�/�8*��_���J݋�2K�%{a���8��v�u�[��`&�/E����\���;u`�e�r(�\�-�(����op�l�{x˪���O��q�,�����x�*[���_��������C�:��()P�^����~�h �>	
��C*�)k,��Z8�l+C����ijIk���k�=@��K�ay�C =P�=nX��2vc����,��@X&u^j�r����"���G�x=���>F�,s�&�����RAC��U�Y����B�%�{��P�D�q#X��g��SN=����u��8q������������y�\Ũ�W�e��U��'��o	@�ii�:���xD:k��[	�<�#��}h�Wx+�-�=?�v�L����(���3�� �hI`��D���?s�F�u������k���{ܔRa���$,�t�}�K�k���ʱ�$A@�V��D��� ����q�.�|jJs-}�����M�K狡���2uO�ߓl�FT) �Qr�6�\��v��� f�C���!���˩%�0��`rKd�I�;���e�����)�,�u#k�q6���w.ϸ(�dp�wR<�v�s� X"���#��Г��� �4�HR?$�[HH
ֲ�*��o.,*I�eV6KO��t��.���ELdU{@�2�i�.$�ԝ��B���t�����=��˨}Vz&u�1�J�Kª~��w8<�E� ���w����E5
1-��E,�bt�OY���۴�lAV`L1�G��X�֏{c��P}�5�hՊXOZ_s��Kql��
�5`s4�9��&���_�j����)��ȃ:�Y�꽪��R� G��G���L��'���Ş]��=N�:�}~�%g��%9=҅�96.s.�E��8��i�E�[�Z����?���7�5���g	c كȡ� ��䀿;�%�S��gR��y;��!��WOY��:�7����\o+NY�����LU���ݫ�_�&���[���c���������N6��TY`�3����
HL8���P��{t,�-��w�-�/����~~N�YO�T�j},eϹ�s��,̋�]�}��7���;���]���P�m�s'H�{#�����1�?bEz�xCrp�ܰ�d=~D�qc�UW��=*�*�s5��/T����m\�x?C��/�a�f���d;��N �x����.	u�n &�DIm�wCɪ�F߸("M�r����~��!�����:��
G-D1�I�r�4�xJ�OH�2�Q�b��ț��[��=q�
$@��^�' av�o��L�+Lw��=��;ob�	#e*"7�����P���]-�*����?�(��2�ÛH��B��X-]}��&dt��$� ���a9$�w����Q���-��`�����H4��~��X;�fߕ���Ͷ�"^kR���m��o'U�%��W�Y�RЛ9�}�:�3ts���mbI��J��N��,���⇉]*>�q_��x�G�3�����̻=�<�f�gÉ�G3����_ �'�E|�ך̜oL�� Xĭ�zE3[.���E0��F��S�ʉ_�	PCX�*�D�\������y�6����)�c�2xKK�ZW�����?��D�����g�g"��G�o�,6��d����.(���:�Dv���z����Q�1n�N��|�¥�p ƌ��]�ݫ��h-�z���wɳm��>[W�w����,��#~=��p�L�sO���9��&Ou-�v�"�_m����MO�+Bz:-�P� 3}Y�t���Fy֝3Ӂd��
s<&���䐲��p�%���=�W��m�1c��LQ�R3�I ��F�\��G�@þS_#Q��Tx ��_DY��`�ϣ�ܯ3�\K����rp��w��ڡ�A��f�B��"��C��NI�����'U�ETӘ�Bȱe-?��Xe\�h����_	�Ӂ��\B�7���a'���T�JFT_�^\��T�/�LK�yJ��k+d����׿�b��w�/�y��Hۦ�-�zh;��%���˽I�0a�β�Zbn����h���O0v��PO�Ǵ�(d���,� �#�,�=&�օgZnUZ7�&#O%0��vHd%|��y�"mC|h<���������l��L��y�-���\���aIr~���$ �6��<���}�f��=���g�Ge&�?&:��:�2Gd�$ �O����.�]��3��U���#ZǢ��K��/N��u�������Yȭز�7���Xb{B��^ƣL9��Y����S��$Pi���ا��� P������{-*����Y�>��6���A�P�x��b�5�u��Z�%A-Kۉ�hSb���&7d�s�.Cz��&E�3s��c{FU�Љ��ӜR����ʅ�嘮^��)��=�C�7���M�p��!��@�B�3�e�S$��������j�z~�뒋&���w�Og��rLty���@�/������0�|��]�d�F_"�@ Քή.~~�##j�w�c��U����W;.����g��t�#I�����H����]a���m���5ɷ�j]�%���r���Xي�aݱ릚*K�y��4=�gT�QZ�z����CQ}@���FA��5��7L
x�M��,Ӌ�}��
��y9�oM�͊[W1�M��Xt J��z�Mb�D�Нb��w�|��+�����[ZM</&��9��K[�ﬕi�k�3�@�<ϟ�������t{�v�� 8ޙ&�&��'.X�E���X�..�,\�������C�RF
���.���JT�����_K��Efa�vn��]�Y&	�<�TP��*��o�2�䚲[ۧ
�4ez2����׎���c��-9ju��.Ksr�n��	��O�X~ֿ�]���5���Q\�_Z<)��C��M�5׎>�������T���\PpMҽ>�, �����n����= �{&�3ms��i���ީ�����P�1>�Y����=�Y3Wa:;7��j�
& � 9��۽��@��0�7e��|�-ߥ4!��z܄�˥G��%&��k]���6Ƈf��9�-ebK㖶D~i�.&��</��.�b�1Eag��^�<����&i=W]���)�z��SC��F*L��9V�CQ��5e��3��^^l�����CB��b2���A��q��Y���hť�3Z3���$Ҋ��EӔm��TKw��G�U[_���h�?< E����OMT�=a�{�ލ4e���Φ�����*��79~'�ɾ�u�uw�"gZ~��g�kVS��y~����J�	�i½�9g�l%�-�]6_��#���24��-&*M�*�~��vrۮ{!�kv�(�V'�t
j�&f	���T�����Jƺ(��20��1_";e#��<��ӶL�̎�$����pՑ�R5���	�˂D���,v�4��Y+eoD�%�?]}�����{�z�<�%n�@��6��_YY��O��6��9�]��He�������f����������~[��_�J�	F�e��ʂ�����u@�{�3�J�T�M<��c����
������.���ELQŎ�W'��F��E�➃���E�ye����ޓ#����ː4k���?��!�>�Cv��.xk�����(k�O�=�7'E��
��8:��mV���0���,��ty.�TX�������ڰ��.Ὧ�z�V3������1�axU%	&�ጴ;:�I��+�q���dv���,���x⃪z��;�xFT���8 JT������ǞQs*�/��q���bh��;��r��k7-hЄ*�}w*
Q�Y�i���\�<�.���{�nk	�G�D�a��y��7��g!Ce��'�׍�2������J`�;,�}�P��.Z�=�����gz�#$P��o�;��^�;z?Ú"�ȉ�����8��j����㘥��,ˋ��{�O��𬋛�n�|����I�w��1K1�����,�{��4�ǧ/)Ws��7��[%����H6��{~�H����6��y�~�$�-%�l+녧�*�j�y�����uܻA6&��<Έn ��Nr~Ì��f��};����-�P��s2�04�0N�V���#e�6��G�ͺ��T�R��@��%5������4� �����$����!ͫ�����	���^7�-֖�������x� Dns�,�Q���[�HF��
_>/X���wR[�,e����t�S�ە)[!���j���<����,v*�8x�?�S^����m��]dRz<�0��-M�xV���}9,7q�~���� �X�!"��y�i��!�[^��'R�KT�N�	��r��%Z��TIyM��7~����e�ۛ���>n��+��5�p������2	a�����-�wN7��x�c��N�J.�|r�>)`M�ů���~i#U�Ej�Xׁ�󹂦�^����<i���E�o8`�2��S��d��O10�r�5��)��2æZo+��DŞ4T�w=��2J��Z��qh"���lJ�6����`�U2��q�Z�nT�ө����-���(O����~�ѧ�u���U�JaM�V�F��]=F��F��8��(7���3��g�K���̴;ߦ�.����L{d�'�R՜k��߹�ۿ���:��ƺ��_/ݤP�~t`�B��ǉ��tغ�9q�[h>yg�����z��L�`�ۿ���xo�~��)��tn�A����~�)a��ӕ��	wC��ߕQ�ǆj3�g��g������rԻ��/�4R���]rG[�{'��`�o�V��w魮��P��}����e���ϳ�*�\�oORW[G/��c?B4_e���]��;����rO+�Y*����DU��O���i���v8��<�\{�w�oFԚ�]����KƪQ(��p�6�@��fi��բ�gR{;�˥ Ih�������wu�������&A�bw[*E?~Ȕ��:�,�����l�ٛ��)7�oc�ﳨ����v*�8a��)�9aI%���?>�(qv?�|[Ԃfάk�aJ�[����~�cN�.�p��j��۫g�N?d.�a��B�*kYL�n6�9�(j5���_(�*MJ�� @w�i����,��Z�C��G��	��H�N�#Dab�g?J�,⯱�������n��ߎ��kԬ�Vq�����y~��U]<�8��qh�m�CQ M�3/(FG/�"�E�����C���޾j��`^���n��.��Eo#�	Zs�����~݁!q%.sG�+�; ��|S��������)��������L/SȒ�zF5{\��{(�i$5sT����ϰ ���F�K�_�t�����y󅦁�b	ϛY�{?��:{Rk�Pl�
x$�P���Pԣ^q۪2($K��d�]���H�"KBrr�Y�(������g�M�h|����&��N?m�����r��Q$���,<t ��dri��j�2H=P�\.���p�F�C��QLa3�*�q�����d��h +�3��^�y�r1l_��V{<�{X�����_�e����b7D�i���J��-�ꎌ_Zyف_�����Ny�"�u�8#J���T�����P���A��m�[��At�i6� 5����hV�>+_��d��TV�ta�3��l�
w�i<;���7В���v�@�lP�ca![������Pԭ�UY���G�9�zF�~�6��w����MCS&�̢ÖC�v��-�
�q��_���a�c���;$u2YP- OA��q^)Y�a���~��/�$F�^*�fNW�Թ��yL��`������gy[�7���b�|DJVwĥ��)����j�Q<MuJ5�l�R#�:%�6���˩ʦy��N��� ���~PL��� ���{qr%V�ty�D��N0י���233�i��7�R4����L���vb�I�Ǌ� �Xی4�=Lq��SZi}$c�'Z�9jc�I%̃g&���΁��tM1�v���RwB~-�xWw���]9��$�l��W���1>|m�r�6$z���c�q��!��m������Lԝ���	�s0�Aj;�
���o7�ĕ ԒGj*8ǵ�Y�xN|ʧ�4�P$ A�?�&Q�S��i�GT�5Zנ���r�h`�3�`�Xڱ�;hm�.��B���������j�U�_���?����SG,��vvz�Y�E7�%~�\�W���*�a��x�%
��=�e�E��˦҇6�Ň�ch����w��+�o�k@d��T�(1�!�F��ơ�����eM�}/�x���)ۧ�}ȣ�4�`�3M�U�Qȷ�̼���/0���e���|��bs�G
�Ozc��cʏ)T$䋕u͜qs�}����8[��nb��ܴ	���⾨���ۻ�l�R�=N���gq�R�o��/���'YrRD&�� �@���>y�4��(u�l�Ѕ�t`%�y��P��@�@
��x5�-\�?�:������>��հ׺G~��z;�_��QM}�]c��C�����������H�tK#%�%�)Jw#� - �HIIw��t	�P�C��9���/��}w��r��gf���~��9��xA��q*~�c�;�nVa#����j�M7^ͺf�3�>�|�)-
��}��#�[���9�)����<c�J����R1Y�rT]fr8ȈI��W��(�=��hHIK[j#��HO̤��������á�����ѹ.��_w�3�ԉ�;E��d�5��qw(�h��4z������_�	;�� 1xG��k=�H��']�G{�ښ_��a�;����֥g@��t!�'�s~Z�&�,/%�;ߘ  �y&�gN����V���3.�
����h�B�V�����{8��a ���&���7��
W��e��k��;}����nJ$����d�x]�z�T���߂�|�����t�Uhc]��#����!BLC���5�b�s��:,n7�b�
8��J��K$��U��G��Y���m��o�ϻ�srp��9��C��=,�1nC��W����aþe߹3g����~�h�������ɛl��O�}�[	x�W%y�4�J�D;hƆ�0�Ϗ ��/�v$����$�����9��贁g�4����v���`�������f1��"��#/�L}�Sax��έ�+KK�m�sk��є�"�N#N��5;�v�
s��szgL�^�(�l�В�}�dlde"P�hl��R����'Y���;m����'{׉S�|��@�3�f�]+V"��l��!�`�ި��-��6��؍�։U;�By�Uc �3Ky���<�w��������W6�M��C+g��w�M��o�����#đ8x�P9"��P�W��L�É��+���Z�����o�#����b$�!S�L�Y㤁:��=�y�dO�N�+�jmqmw�r�� ���r���V=3`)�ؤ�3S�e\�X���,k<=�+��
\HMD���^nx��ާ����gO�p��D��h,�?x	�-�O�(ӭ��Fl�<�Ck�e>�Eg_	��e�S,�E>g��D�
*��[����pEy%�JG~�
*�2L%��;ڟ� V�CgFd���l�Z�>�c�&��-�T����8�T�$;�(иs��Q���7KK�[��h�M�{�
�hl��!z/��.���2��Vtfn��IC( 3�,͛������O^��n$�c6�� *6���������U��k��r�#rک>J�]�>�����b%�yK++0O�x�C�;��S;�6 v��|�J�?H̿o�x>���mi��q<{�;1+<K�"Z������^:-�q;|1+���j�����+����\C�dGQ��Uζ��ӵ�<�ZN>�$��og��"�~ڋ&��Jc�y�g�g���
�L����ʰc�{�7'��-Խ:S�:F�C�%���V�o8.n�5$v7�uZL�3������k�����8�|��733������tW���P�%)(��o���Zʒ�λ��ٌt[m���n�=�ZW��10�&R�Y}�a�jA��Ӹ�0�1y~�N�
�۰o~ ֧1��=����@�!"c���mc����G�.����Kg)���鬮���&A�Xs�R��f�O�s@[�4����wh�_�ȴ�uձf
P�H��(J���z�f�k$(����<8<��Y98� �6�\����c���	C��C���!���i��_�"~�%py��s@�[��G��
�}����8����'�u�O�(
]&��`��h[��+�;��uO ��DD���H.��w�"5=�
P���؜���e:��K�\U0C�.'�F21&ڠ�Jw3lf�ݦ��:e�N�������D8S��;���D�(m��@����xؚ(��\���#s@�͍�DK7���N#^�B���H XA*�ٗ0����%�������� '3�	4������� DX���#��7�W� Z��Y[N�I}/��u<�E	3�Wk���|�Qic�Lx�B,Kt�2N�]����`K�쿹)80D6 Wz��Z����;�����h�Fɴ�Ƿꞔ��LU�E���Ȕ1`���2@�[�����s����vfV�����u�`b>deQx/1�0��P�Qh'�-��,\6��/�텓�LC�j��Y� ��	�yW=�hϗE+��1RRR����s��e�z����%RG m���Y�6"�h��%�w����jq`` ��=����.�]�����1dLҸPaξi�d�<R|#?��C� J}�'%��[S�̺5z����yMؓQ��2��kdf*����M,�[n�w��!h5Ba��,Y�n~���EӬϹ�Ҿ;]g�9g�>`D&d�|l�B����Gd�W"�;V���OSӸޥ[Ih"9�]c���@QFk����W���t����9{N"�=i�q~���/-a���t)���[��� ������V���w�������I䂹��*��'!*������;(��U�Yz[8�'�#j5�K���Oc�ܹs���-C�[������f�}%�a���D{�=qő��L����A��L6�Q�Qb:rcI�#;��Ye�sq�==��7;��ҷc����_�d�:�id�,�1z9�e�9���!������r�K��N�ʐֆ}Q���s��m�OG���!��;l/oo�������� b�rP��=ز��U:5�P_V���� ���Z��$�y��"@*��P�͝�ƀ�f#�v�׀��������˧��GT�+�r��zL׮9W��Jf�ѭ�[��y�	=9�z�EJ�J�g���jz}�E˘؋���O
D��<�*�o*����-����Kl1�w��nNHA^�i����獭#���{�d3�tI�om�
�nYmMU?h ����W찈�:�%H�E��7CԐ�]�@�X���@GC[�Q��Қ���������R����p�>���֑��h�e-��,^t:R���
�%~H�����I1O������zQ������_��{��ť��פ��[�bF�K��:k�|!{0N�yW�� ��_3Ύj��2�U�W�ˍ�ww2P=ަ ƒՍ��Yk����H�هd�k��}]p�QeIDu�R���������$!!IIJ��������ZH��>o$�n�4�ΨaMFH8��$��!��k�㓮�ׁ��9[7���Ҋ"@`��&Pz�r"�=ߨͥGRן4�����M�V_
kk5��X��<}-B�\����K0�`��tO��c��T��a^x�W���]�r0eUF��O6fye���� L:!���Jˇ
0�yW��7�C��UKݗ]�\#����z�6�]aR9��f��C-��q=��2g�Z^vEƗ��<�����~6744��n8ZT��0w�䞞��1;���v�P��ǳx����Aن��������ihm�[��C4�!pf���r��Ƹ���;%����@;[?)�������l�D�gz��e�Z$�� ����d�Jr^!@L��ƛk��˔<�,�5�	���+岦�a^�kѣ� [�1��P�Js��1��"2 �WqR��`��̟�e`��ow$�΂c i22nf�I�~=P���4�2�z�~*(wdo�������&��J��D(�\?|��A��S��jA���{

����A��.�ߓ3��lc��8��������=$TB<6�!����A먶����x���4DGGǘ�NQ="�G5�#�9ZL���@���°�#TTTB��^o\�u���R ��Ϝ5/0Ho��lN�}���v
�4�1춎>��@l�%�7���/��R4/%�ۥFVx-��qN����ùh`_@AA �cI�B�	DP5��U��+C�xg�R�$ײS�¯l
h%�*� �ڐ4�� ��6&���ނK��Gn�����<o	f����qU���=pam\/��e\�/[x-�VĜ_/���� �MO��<�].�q�p6
�Ӈ��9p>vZ��N0" 20�G� ��~�Qw��p;WL�b>H>���_�6=ƪ]�$Ϟ�#��Vh�Aܪ#�%�8<~Kt�,�t7���夤��&0��Jp��}&�x
��P�ܥ�v��f���*��0�F����yˬ׾���ӷ��j A�ٳG��=�!�\ 	�r�:�icIc+��9�~q�t�kp!�3!H O�O��7�}%���?�����6{\�ϕ�mbd�x����2�N��4�`���^�ƣ�y��<�A��A�G���2]ƙq�q*��OX�i`���Q���/e57$����
�7��GGG�j�'���MsU齏��6�ZK1}O:tZ}�?d�
l�D
��r�|��G2$/4O�
��O��#/�2���MMiT2�������0�@42�b�8���r���֮�0���|lb�Qo��ف���nG�V��5��H__;�x��Ӗ��D��O3ė����>�&��T�\�|����t�taB��7N�ԓ���nٱ26�XXX��}<<<�[�v��^�Fؚ����7�m��~9l(����"5�)hg��.�G�Z[�0ܾq���c�p��ȍ�;o�i
�yy�\j��"�~���ҽ���f5����Lz�e��Wz�O[�vD���d�8��~�ꒃ��q

꯱A�d��8��3` #��TٓGݏ���*�B?�d���2w�ϥ��nb����bn���[Pyp����~`��@�ǟ�Q�8�яQd���n''���������<��;����#�BDܲ���uZ?�88rV2|�#�����yy�� bC6��Ah�Q7˄�bE�����9�Lש����|�n���M5U�C�+zxx(�󰡱��r��(��[E����S�?�p��fJ���Gvw?�9�JK��:�z@��I�����;^��٫!���Jd�&-Lman�T\\jn�����êh�)y^s� ��^[���YÅX����zY[���+�yGtӫWZ��œ�R�	\������8~x�
���e�Օ��������/�+Q�Z۱tAO��F6�56�t��I^%�\�Iڃ%y���D��h*i���}�.�e����PSC���:���=dz Q6����*� tK���s>���HR���@M��N;��c`%j:�c���Xnƈ�>����#��z--�I��� �;��*b��2�'�#�R$��-����������x�]�
�1��+��>[��m>�-�߮�9p����h�-�ڭ��,�FW���d྄�&���i�P�b���(�����̻P��7$)6��>c�� ��@=�e��U���� v���,|��ݴ��5��x�šP��[���aK���
��!��^���c�>Jb��CK�
шߔ���H��î7��bM��� ]���ͤR���w��V��s�����:�������+�_/����-���� ����"��=�-d�A���P1��~���Gl�7���6�xg����/�`A���H����ɱ��ފE�H� A�=m�ݰ��Rp�&�UcS_�8���nЖ�n9��au�m�!�k .^�����_J���QVUN�1
.<vh7�o���Es�WYѥ��@y,� �a�E�'9`$)�O[ʀ��ή�[�@O��=�U����^`Ą�8T�uЕ��|uO��ؚk5�k9���V^^TL*'e#��a�5���Apǿ	�Oa��������5!^ޤ��">���t�t�pxo�A��3nV@ՠw�FF�x�%��;�u����Of���11����������2�7�GQ�d�G�C��U������+T��|�+/^����XZX@G/�N�6���	�.�z,'���:��EJ�7����$�z,��BC�A8<?���K3pH�9O�Ș��#	 �T�����Pۼ�VU`֘n��SeR<��ص좏zL�����������2���daz:�21@2Y��a�. pF���ƝsG��&�z߄��<NKC-����?k�^^M���M`J8�<��C_�M}?Z���+D:7�!�<����)ͱ�|C)�G\� Q�ߨa5^m���=M6� 2�c���rr��K	�_�{���;Y[�)ݶt�fYZ����gC	@'[9;4�4�� C�xyy�d�ͅ�Y������j��&B�r�:�%}�A�)��bG���R��/]RR����cL�jgg7�e~cֹ�J"v��J�Jچ�߼��V'H	�Ywi &G
�����'���e���y-���0(��wa�4�%���q��/4�8x��(HlO��7��#P�����s܋H��y��&���b�k�T�{%e�ӵ��M�sw�&��,��Ӕr��ąn]$ ,��ĵ}������R�ٳg�L+��п=F��-����n(@u�������d���]�ѸE�⩇��=�>���2@�Th�x�� ��:I��RF��,�X;���2�n;Pr%���.��wQ�.ll���J#j��)����y
,T��R:�?^��/�4 q s=@����%(Xbs��E"?���V��9Z�Fu�����Y�3��9�ctK/G!(���3��he�𒖖���#��׻tt^��ns���]Vb��T����KD,���ܪnn��C%��J7,��~��I�������2��ƿFio�X�V��oK�L�l&y�����C���g&��xy݇vD������i�l�A�&Z�2~,���� ����P����񳖺�^bku+���_9�VP�|$�-m����>��M�ޯ5㸍�f	��䏛�nF�}�)/@ό�E���$$$�VV�6�4��ٵuff����m��P��m=;;�r��1��,���ЧC)������Ȥ�� C�]�������Jo������&{2��Vxxx�)=,/��8%�IO����k�ptMeL}��f�gK�?Sq#���4�������§y%�hN66����ԣ�>O�꠴��ܳ�ć��s���g�`�lo�܌�pu�����s�<Z�-�V̇P��`��|����weeZ�i��q��g�^���B-S�,L��3i�_����#N\Pb�˖����	(��8��_~����*�,c�6)J���p��� �1�y�gg��3�ffߝ~��������؜:�������22XI�?y��j���ۍ���ө wX=�3�'`�GS�*��!	`���#��&�B��c���)�Ig�N�?(|��|�U&��,�} ��)���w�@߁b��@�X_[JᲒ�����?�*��h���9:��{�uq+�{r���>Q����BzE��������^���\U��@_�����n������{�M���y5j��8�+P�Q������@� �<��g�d1x$P�$���=xP0(��)�B_����VQ*���&
��榚��{]ݱ��Қ��ax��w�;G��"��^hm�ƫ��4u���y8=.�,m,�2_�������*���[Q��w�\��P�����VNBD���� �2Kn��]��_��U��>�F����6�E��p��i�e�EJX���|aikz����Ďì�{2ǃ��W��O�kk�����^�)(( ^Vur�|Q�P����� r��4��7cv��]�4E�?��&h�aL쥏�^3ζ�!�ݛ�m=\���Pu�qY����xJ �*�<V�N��E����HEق��f��$�{��\q+!_����*�*�����(�Rr��g�zJ�#��#�$$͋�:	��K�T�O-hN�9�nn�&^SEw#�ofdy	���
��ڝz�t��nL>X�O�E�i���6S�~���1�i��Nrڨ˹E&Ũ�_� ߀K�j�����a�<��_�6y�[bE-�!��K���*-9򂂗�B�{�τ@�����uK����\27�߷���:�2��PHH�6���S��־����G�������P�=K8���7)�����O�^Q[�ݟpI���k$HЬ�ڲ4��F�8Y>M�A���Q3��K�à���6����K���� ���%�� ����g-{����'��)��-X��3��)�W��߽>9��^�Oo����މM���z��q+<K0�9��7����3�^ٍp�0w�*���{F.��ι������ﾃ��� �/�d�c
h'ܐ̵�����s�S`��5��twx~����0M��c����!he^Fu��P.��G�ed�.� �o��r��Pu(eV$��g���4˵�ʵ�">W0A�cxxg��Qu�_��0sr���;��L�E&�b�?5IFD�-��]x��"rI�e�L�����겇���!�\�T7���HNo��o'�b>�APD��x�'������C
��w����O2M0���O�����b�2��Xߵ� ��F ��� ˈ^�퇍���LR&�[)h"c�p�l�:��5����K��ؗ$^���R�׬4`vh�� �z)"cpZ�{�T�\˺3l���
�(��X,B��o7p���7E,ۀd�e�Gl�X�M�Đ�A\nB��a�d���4����I{S�`C��]���(&kJ�y��-��Jk�����,DQ���Z�--��w���h��H���,Ӄ Rl�ЂG��6�³ #����Ng��axI��Z���N3�n����#	��F�8b����\�p���E:(o.*V��L��t��G�
}��zG���i )�A�W7=�r�0h�H�k`�x�噥"YO_�[ )d�۔n�(��S9"�ɁLhY�fYM���9��<jʔ�>g��/��˦>��'�U�K�d�S�\�8�ʰ~.-%�D���!���\=���[ )���
�����^��>�����v�?�tz��8j�Yv�id4��*oʃ���?����s�[���2xJ�/�P*�����θy�͌�]X���������;ؒ��6%jŘ�p׵Z��|�:�9���=h��'o���������κE�l������TU6.f����^щr=�ˋx�&I	�y	x�fR8/J��{�k�5��Jì�C�#��IVƔ���w��%�bc��
y�K�fӂ��I�[��ٓ�+ʌ�dnQ0��T���� ~n]��y͸f�]b�F��nuuI�e�8K͸>6#��]~jc*���c��92l����﹎w���I��&�ȯ�����n��,�E1��k{F�))� A���K?��,�PJ>��.��Q�����&@U;9��y`������1�gx.�[���ǺR���-]qz���ԁ��ԙ�欪�P��C�N�L�]���]
B޴qAte�T�XҺ��c�CN�t�&����Ƶ0����:������g���ɂ���8�E����T�j�*=�u;�R+9$$HΕ@0��+�HH�IB���Թ֚����@�c�/2�_}O�^�s:${���h(^Bۇ����||N���� �Y�ԯ��Ȝ�I�;��_�%w7잒�}�z8�?�'DE�+_,+j��2%��Q�s���Z�j��-�C�:&��ȱ��.��5J-�in��ʢ�)�'�w����P�X��R�	�}zd�Uզ�5>���+�Vѻ�c�x��;e�˼Lr�G%�,�Aᳬ�ni-���������j珘n����=1>D�{R%�4f�1�5��K�ϳj�v��|RE��Û�lB�tsS�y����j�����W.���/6��cN���Y�GK�E�;f�i�/#B6]����n������v��Q	�ѿ}�"��l}��6��A�P��H��ZJs��H�V_���l$^-��?��X��W��t�|w@�75�nFV��ωԛg|�j�`@Q$��%,&=$l$t�����S�(��u�`4]d�&�'d�G�o����q�?>�
��_TSx��g��:��=�mRp1����^D�U*����_�ñ�oM}����ΆQ6��2�����}� C0�+o�r�}NG��4m=}ve�^R����w�w�v��o}�����i����Y�X�MJ�Y;1P8��EJ���c�jsN�5���eNB�ߌm0|+�ۻ$������8�͓�?�N׻��\� �L�;��0�c���,��(�S��p|�ʜ���5`{DR��2��kԜsвZ�!~p͙t���N����'M���-'?��jrz\���D��6�����Q�����%>�]~nl$ZMM���ڹ�Th��1���p%	"�V=V���=
�,��e��0?����_~ԗ+lp�ʴ�O�O:%���Йoz�C������g��HG��)f?OuĦ4-�X63"�$� h�?!]���^�HM�FQ�m��׈e����/,`��D���KHJR��J�`�	@�]ZR��o����xz����������IvV�i��D�[����s��m�{ٴh��\!ݺ袹s�Cn��Um�sL�����+ � .//_!e�!@��&8�Ü3]w�C�ϣ43��H ����N�KHD���^ZZ�r�e���|��Q�oT���(ŅWI��kX,a&T,���&�W>�9�~�V�|�-�=44.nm�4??���rWBJ�9���5?h˴���֖���(�k��DDD��u�&�𖉡��T���*Nܟ���N�\1�<I����"����q-�r�N��p��5�;�ql2J�[O���UU�����~� 9P�%Y)g�\H�too���D��o����Nd\\\�<��B��;R�t͡�u����}�~I���z�KP|씠d(�aƚ���#$*̒�v��C^%�޴�V�q�]���9CwaI<���Q�W�X��eV77%@l����w����t�����#��8ݟ���L� �o�K^��|I	��m���6"s�>��.!�M����fRhh��R��(���x�Q��;�?n{�����p �Zfyl|<;/�N||��u����j��"�/z�*��}�)��ەr�Ya;�!JF����Y�1�Z�]��iM|�p[T�ٙ3&&�]zz$*>9;�#n�G�A��������������Ȋ
���Ĝ�\��].�^�웟.���Tb5^�a�B˥��F����{��|�Pי��ꇉ�
ntj��P�G�TT�`� KX�ß{xxd�Y"�>I��,��M}ਯ�oEHGG�+��72P�F��(F�.�/3���QZ�aqͲ������J�wd��ۜ�R|�V>���wycccr

�����%��)s�+M��ss�@��>�W~�Q;�E��H�.�e3������r�:�q��ylE�ō#ﰣ3>�A��D��*N�4���{ڄ:�ث�U�RR�===`>��r`ή���{<Zi̙���ܛ��EFb�
�����&=س>�����Tޟ�a��U�`&h�Xr6LI"*�y����Z�s�]���F���Opg�UL��C+�?�N��:��+|�q��$�"alL�<�u�"s?��{Cè��;���hWa��C�����>6���ڊ]��(w}�8��du�7�fV�O|Jg!g���qtt|����iF��Q�:,4TT^�t �I����^���M1] tyyY����Vl�S){���QRl�h��b|iz��Y�t��d�C|���1u�.=9[�Q��{���8,|���}�\4F�")!�|g�9I���)r\w����1����z
ۇr�V)�451-(N�Ho��e�kb%��K���DO�-Ĝ�xLz��׈���SE�����&����5F��j�u=������`"	&���9�f���rr����3��M��M�<��e��o~��>�� ���~�E�w�	s������+vVY��KN~��_���wqᵸ���:��;���q񮬬,��0R���C�|� >�y��r9; |7�Vo��$S$I�LPK�T�5�k-�� v��!���9@/��1�x.HsKK�g��M��jk����,,�2����3̼x�)����ɘ��d��N���m/�,����@�a���rww��Z��R���ۏ���g|�~�6���H�b����� �����[���8|�χq�J�|���S�s	<=����T�Y�dR�((���[ɥ�n��fgf�F򕤍�?<xv'1)��ɰ��7�����
6
*����C�J|���ũ`�k��W1-G�Qz!Yśaˡ�����Ŋ���K�̽���U�g>�������S��Z��_2���m�@�k���	cv��
��Ǡn+�����,.��?����>�mT9����2<İ=��;ra�jkr�wH�DK���ˀ�(���or<6�'^\\ɺ{U��4�Mz:)(ٞK'|i��
�?�����?;XM�id<�3����~����~k;�s�Se��λ���`t44H��$��$;;�)��H!&�\�DI++F(<ZZ!�|���&��{���M���{�bI���~�f�vv�j;�T��G���5�_�C�n]��to���$�l���_⣐��V��1�Z�Wg�����G��ض��U*o���
�����oj�Ѕ.�m�k1g�M�ؖ\hT"w�<ƪ�xr�!"J'B�,{y�8�q>\t�l�Kh������1����Hb��j�s�±u�9�bFe=��55���T�$�W&��e3S�{r�5��a+�����N	>@T�t�Stl�B�s3�h�z��X�﫩��Q�42��t�l=��t�^t��k��I��p�,����}�G_)��(b(�Ia�����+�+�iʞf5�&�� ���+ʅ�?Q�v��سS>>&k��|�~�M�Bmmm�P<�Vv���H�we��L'��~���s�W܊B�?�S�"
|�l�İ4���Ո(x�$���e�aw;m훰��������h̚��'���EH�����>ɗ/�"Ʉ#����\v
��KW��:BR�g�CC����F//��/P�1KOcb��z_�k��)�q���R03�k�9 m����ݲ�˯W.*���3� ��B�+�z4/`C^����}� Gh��Ej����ݓ�i�?,x�����)���D"���£�?B�Ȉ�H)����e)P��|�w�d���J��i�GB�����D���4:&&�Ouk�#saA�d��y]ؼ���(�5A��-W�����宮���p֯��Nb-��zz�� _�]]T@Q:��w��>r�8q�a]�r<�&�������P����`��+)���p��� �4'
o�������r�SG���
ç�|$	,�a4r	�uu�n�_@��8޷�iL3�=%�:j
{S='��N��PHQA�@���6���?i��������'�~��D����~K�fR�ؓ�%&C� K��\�h`���P�l�ԛ����b���P�or�G���	�̬�y�H��U���s�+!�gӾS7�9�J~n����%:::?�0�����܁h��t����G(O�}���hr4���N�q�N+����u9
r�N3���kp^l��^o`?���.K�Uc`s��+֩FED���k�ۀ-�=B{��|l���O�6p�PB+�	���I���=�GEy��<b��x��T��$��^� �!v�Y��iA�ѫCQN�]�n�	?�����6S��I��Y�-�������;ý}�E��Ǳ*��c5Q�Y�߸ێL�V'� =����5�"���`>���Ob�9]��\>�,*Z�ɗO��cm�]�:�kSQW�S^:��Sc�~�>`*�Çے�����G�	��9{�z��Y�BM�Dw��9t=��s�_�!"C��a?�i��D���ZB�k�i���R�}�m�����J�Ԅ��5��[���$0����~G\�e8���0�(1��R�0��쑉K��> n(f��}�=g����CC������-�r��������;,̍Đ"1���?�r�)_�r젓�����~m�׋�Ť�e�	�1H����~�òCRS��S8�uE�u� �{7�m��oT�\I�;!F�Y>�aV��ĝ��`���问�Ej���5{h�b��5��%%�0��@G��(���{}���S:��'~�͎b-,��UL��}�Y��_���n�����?̼��J�!~�!
��DV(�л��\�;|���"��(�����nZZ��i���H�YzYʐ�z�*��'NBt �?�Q���n:�}c�_��~��ƌ9��޾�Ty����Q�y��=��<�o�]�
xhP�O�oC=tϗ�~N����/.�CBC�T>����~߷�X�L$��"zNNN�Q�,N8:B���|o�X_��ج:Ռ�U�^�tP��Jďϱ݊�t��K�R�
������	�ne���x	��R�үY����2Z�lht����� �ɽ�
AHC���*�(0Y+Jo�!u2�0>�_J�a<(�͛5,�	%���.���;ctg>$A�'��UnZ^齆1iOt���Asp��K��q,�`�����T�m�{}j�)̜`L�f���-�=n��n7�.���j�֏��*�����9��
�YrA� ��֣�}��}�����]�8?����c�/��%O��#;�1��k�gt?!�`�EP�k�g$��f$9���h����'S-A�N˷�ẑ����Q���r��3K&''O.�T���ܳ�r�W�V���w?��&��k;H��67������M�Л�o�wo�t�p�NV����i�{NL�`�S�D�fa�s���k���^�,'��v���M��uT��HJ��L��ۙv	�P��𯫜����n!��Bmj$pB�O��鲛�����^��� �UwyWQU���sqq!]�o�;���A���ХCR��%0�Eu�>�^�;�6��HS�H�7���S�e|r�����s� �
JK�n�4���5��������z�����=�o;�,�*C���+��'���>�@�y�E6ѳ�b������^�o�i�{���-YW�˼9{6,��բ���4n�<�	����a�w�P^ٜH���v���w	-spq���g��Rt����x.
����bï�������H�Z��S�f��gcHoƘ�?GNM���r�>!Y�R���]{�.�������d�Q��ɀ����U+��u���oAÔ����1s[�ga�p��;��?)3���(X#�E�Xb�52��r��'T���T*6����v�#ԼΣw+^T�ߑ�o��N)��Y:��r|D�����*䴟�(}4l@����p�$����Y�Le:�$�ņ��_�<�E�$4�t�(���0���X����*ue��K����R���#���W$�V��<����tku������x�-�^H����Cl�\+W�h�ɝ@�G�uk*h���;x��=U��z��+,���-#g���\�J��{{zځ����Y�1^�u�n�+Q��/���߽斖�y�l�6VKOn-�6�}�s�J�	�7�M�����k�wK����Iv+"�������=t���-7at���d�%W�]TԎ����c�_���m̵��ב�o���օy>۽-�[z���֩i�z}\IH�`
���n����#�α5Q��`=�n;X�8�Ǳ���|/,����s���A�r�	ޠ|Z�W�j�1~�!��f�M�vC��5к@��[�1�d���O�WZX�|�����;52�_wH���CS�o�S�5 ����|a!��Hr�w�>�
���u䷕4-�v0l�\���~sNª��O\򧧧I��<����:��8knw��H-o��S��G��wO,i�m"<�>�s�/#+�y��}tz�v�s�/K��{�񲸸���� a�f��lc��ϵ�|���cy��q�F@L�J+��!�(��>����B��P�S���`�̬����%�C9����Ƴg�pϞ
S�d?��u쎇�5�6R�����*������� /qpۍ�- �Xئc�Y��A��e�JјV�+6v��\P��1j����`bv)pϼy�a�s)��Hk�Y{J��R.�k	3�n�`������f�zL�x|\'���&�\� �f�ߠ��-�)�N��A�~�kVC����'I�o.���Ѝ���79E���Lq�ǁ 7�ֱ����_86bGQ�����|o��
��u�w��B����9��JF�����8	\�oD����
Z�F�f｟Y�!���a�L{���e�7�,?HX|����}�B"o��*뢐�Hhϡ���˗`ʃ��Shc�uvvv����e&ddD�}�&p}�O�̼��"g-�h};"߯I��>����!238}B8w���$O�c[��q=�=�Q�2�tJ(��Mȁ�H���V�Һ��1�XDh	@�ORv�?�`"	*�e���+���-�G����#��
�E7X�Ơ���-}x�I:��&�����	^� �ң���]Lȭ48s�L�ߊ@H��p��= �\1��sQ�	��V)�/Q�U�i����BDW���.T�]6�EW��"��~#��4/����k�wy��wZL@�hs<''�u��n-C�20 /����}X�q��)��bf���>*`�r��9s-��_8K�]x��Y}�Y<((�d^X�ؑv���6`��]���4�sK�uZ�L���9��u0�@�EAJ`��w�_�?.�1�����*��[:�s-$R9C��)<{?��5Iw�H~9�Ld�t���u9���܎n����VR�R>Pz�һEo���s_��^wSt�|��pͤU�y����.$2.rrWy4Z��� ������ZQ?��������d��[�v�U��w~Y��ꞷ�ͽo,�f�?ź��'x�����?j���(Qq��bO�G�$��j���3M��yw�~���i-������)�(��,h9�E|�L?���P��zd O�*~��齅�K�.�F8��8t��e�PX'����d�T�)�����gi>�v�/��C��jU[���Π�)�8(�g'����))J��%L��K�
ls>�e�{��4Ү���r��;_:;Oy��W=6�slba=Ɵ��N�W<��@A D3t0T���|�/�%*��9n��C+��}<���uΣm_TX���Ə"��E/��l������C���g��B{l�WύZ�ba����� T]��C����48��Α�eϲ�"wsG1c2�t�?���J�K���Ç�3.��B+�FFFEE�no�e�o
�k�ó�邳KhK��4�'�<*G'&���HV�:,~�M	�7Q�H���	z��}}�ax��j���,���
�-��؇e6;V<�ݖu%$�]�*_�Љ�/'�ϫ8�����g=�W�g�B��X%�fd�Q� 
��������V��k�s�@�k5{p�ZVc�"a䪆��<�z�����HX���д<p|��D��U���_�[�q���=?�
�6JĲv�~�����1�m�� ��\-`�^n]{����z먪��_���8t�N��D���;�	E��� ���%�������{���d8{�91�\k�H��d�6SR�;'ȅ��P�5?���/"�t�+��eRg��]o�g:��Qi���;d((��R}�c՞gf�s��/��F��ӷvv6W�c������ζ�nj��	�]�i��h(�xS�'�	�����z<���"f���rbb�q��㢌���t�A�M)}}��"cc�S����6-��#"m*[�)��/oz,�e Qc"~�O����h�^���Dn"��+ �O<T���100|3X�������
�^���x����EYpa����Rr�l�\A��<���l��j���a,�(�"�t��ܟn�$4,��Ċ**G�0�腋�dߊ�����at�ׯ_�r�᎑{(����a��i+e���ݍwFB�V����]�w��8� ��EԋU^���n�� ���a�O^�qb8u]�����\���'�N�+v�H��mfL|�����n�;s0aO���Z�D;c�k�����d���'��q�j������r�8w�%/���r����P�J1����g߿��O��z�Ժ��'vc�w�@7�qǭu��ohh�a����	����������PI��t��%�������]ZIC?�MQ�9Q�|�}#<����>j������q���� �_n_O�iVW��:�?ߗ%���$\r���|���$%�)��/r��)�`�w��#4�ū,�~��@�)k# �����wm<�hN��y۩���so���䎌�J|h��z_�xq�|�O����H,
x�W�J�����סEC�_���jk\mr���ui�����W�}�.�Հ,dL7@����-z�@hA=������_��_^�,ں��o~0nxF����;���+Qh))�Z'i,^W\ ��R.Z��ԕ%�|"a�KD�� ����I�r��/0Ub�p`&�s�/үa�����U�ݨ�`�h�~��=$id��K��X 8c)�FW5���;�:��T+lll���ݎh��oF�p&#J�)�unl�y;����!.N�����2�q��=WQ �Y9�1��P$O��U���
�������zw���;�ߜ���<�X���� /l��#'ߥF'�j3d��+r����@�J;;;�c.D�+}��Z�Ϝ� ��'��<��,�[J�K4����S����6$څB���r�����y�9��Cw��y��*wQ���4.phZ�}��4��|�j�o�,|�9_h�0Z��fМ0Z5��-��9O�.��M��}P�*��RS��ø�5;����X�>���$�nc��+�~w�4LF��o�B�=�4˦a���!�%�٢�iNwB2�1���(�H�-Y�'�\���r���`��/19����Du�K����.r�?8�Cb(�<ɶ +	 ���p��u��X�W��ͧhK����������|���-)>~PE��i'j��ye��������u��m��|1u��;������i)�׈/�}�x��6���6��Y덏���������*�P��QI{;�L&=��0�ri3��T~42Z��^KIn��.M��/e��9=j�*�C4���ɝ�X���ӵ��f��8��}=�7���2D\��lm/-Q��F� ����߾�HH!��5'e�R���Ӻ�^ڢ��y�kg���rsss]{9� vi�|����-HJx��#t�R��(ȱR���+��KGo����~�ohV�d}�9ө����IJP��llN�[�aS������jj��;�a��:C���عM.l%.R3?���>�u�Y�h .=l���8O��e�Y(&��5�g�~��	%�U����,�o���IͶ�kE�Ԓ�� o�^��"��`0�X'!��[�П,x�*�id����2���܅p��G���ߨJ��!�p�[�hO��}.jv��Ƈ,n;��#<+��f2;1_2�����	�N�pb��(L������}Y�m�f? 1��V��1�n),�w�WH&�98�1��L
�A55�c:/������^��;> �����<v��@�ߗ5{��1�؁�|Ř$jQ�ޠ�D�G��!����3)��
��lQq*Q���G��h�;{��d:�̈�3���3��s5V��z�(��*�TTS�;jX�/�������L�Y�[px6Ľ>��Ո_�A��d�JBW'�@�_�������D����]vE�ϾO�A`�P���������	���a��d��MŴ��*P�yQ��|��)���Eڧs�P�m�K��}�M���n�B��(LL�
����~G(A�3u�F��NN��?=u<��A�!�|s"	1qx�IE��HOOo���]0������>7�ٲ���Ѯuu���*/j���k�Ȯm5Cd}�׹<٪v��tLL��ғ�gֱ�)����T���TWPZZ:�ĺ(�\�:$W�����)#����A�{���:�_�(��)[�#Z����Omzz{�s�*0��9~�� $HW(:AbN���9�3�Ъ/��ぱ�����0�x����\�H��.��b֑[�%�h��*��/��W
aHt�p����5�> �L̛�����Gǹ.QuW��<Q���պ�O$V����q��n��]�JG���ŗ���"��T��A���BF�7����ҡ�"�HOn�\�j	D)�i~�0ڰ��r���9��w��[��t��/V�fN's���Z�zO#?�U���g%���N���� ��
Q��KCӯ��Zw��������S���K�^yo��J�Ԕ��7��"#מ�t&[��!�+�����_[��Tr�r0����0�Z�Q��g����S��0h��0{R��`�����۷�r$R�E4o2��`�F--����-�(q��'K`�2��a���v�n�җ�P%wO������EO�� �zG�lv�;��d��/�x.V���-��Z���RY�p�ka�BT:���KZ��� F�<�%Rs��U�Ȼ���F["Bm�����|���Pv�;� fL�`�NBd^B���Ng�h��ѥ���	qT�¿�
�����p%d*~��W�e�X����ETT���z#�2��y�¶D=Ry:M�i������ܗj�Ҥ�/i��bTf-NO#�� [,�\?��������\�B�4G-���ѐ� ��O#�K�����̃����ZWY�9`� ����e#���A싧
��=�w�ݪ�7�;8��6�a;t�$K�%u)���lؖ�Y4����ǿ)�s�̓�E��[�sttt�qL�x� B��+'���.��S����'f��#s���g�YL�
'q{{ۯ���a(�5��H�Vm犺�q��n�|��^�����rH�b�z��l�u ����,��$e͵��~�]��m}���|���ɇ��x�	䰄ҳ��3t�nn�pm:�6v(P�
�І3�[7���Y�o|�e�����P�+N�� g��A��*�Vu(�b�A��hBZq(����}EH"o�G:tG>m���j��6�� ����I�����w�I %niJ���=f�t4��
d���$$!���d5�GA�n��"�Һ��M/FG��/�V�D7���:�4Ti�VP��^GwW6����F��"��+�c<lU@^�2���%��\�?�gY�4t�qeєg���=���c#@;��沐Ϗu�B�N��Pq�ũ��]�0�3���AߵX�ߗ��[GGU_�<e�������0��`���ޫ.ّ&����ַ)CP|�罴��XF�1�2d�Ǐ���T���,�L��jg<2��)�I%|Æ"�����!$����H��F�H�[��mXf+�h�b�s:�%����x��1@�N���(<8�۾�������U��0@��A�Z�:���
�q�I=�繁�����'��U;��u�)��������<~s�000�ؼ���;�u�����Z����w�ҺX&�YwVu!P}�2kl^��ɕ��6p
�yV��e{��8R��0�v3�
���d�͏��F�ER�Py�R�to6q�8��{��L��;��Yב��ʊ�����*<��~6���5���+�Z��Ax� @��Fv���\\�
	�G.=�!jx5{�h��jLC��S����$[]�����Z~���8����;���ިYe�)���e2�fA@}�Y���3,�_�ˁ �G�V�O:��r�o�v���ػc�fP��X��D�h�6���E�ѯ�tL�E�4S���7�8�E�F*��K��q/�����3J�T��8��H0�Fbe���FvbL���o�����߾�J�����Ǆ�_x�O�t�|(?\0����\N��l�+�tc|;��Zf�,~�΅���zn�cs����8$����/��v�h�X����H��"���9��f| ��8K��.�u�*�K�g�PV������Fb`�}!�a�fKvtry��F	���l���144��di{$�TK}�2�'��=����B��0���6,p�g>��KGk�f`�R'u�X-��x�>}�*H)��~��!�w7i�����O?����=k*�0�� ��d87���h<�܆F@�6+�up�R�v��0�‎:�	�m��o'��f8�qF	��l_y4>�꽂�t���o�F�Uqa�U6#3<����UGͅ�ƿ��������p�)����Փezz��o�c��~����N�OI^�!8��8ݜ������F47c'MrQ��W�{�_�`,9qg���g���V��Q:w1N������W#0�FFF��m����3��F#�G9��*
 ъհ�uXay�L�Y��s���$S����n�dz��O�aSl��	�}�m7f/���' �,�����w�TY����Ĵ�p��k���	�i��LR��n:}i��s�o�D�d�*�{R�c��O֖蚶��M��Q�͎��D���� $�g)G�~�������{�B��o�~��W��Zl3#q$�Ja24�0�Aa�!R�c�<"���S �*�P-��C��Y��b�V�J%����%�Gb�I���S���/�){#jI����}(3l�+���bR301�����;WOV�NJMOg``�^���r����p����C�я�j᜖�y	���UBi����L�W���qs����3)��M�A�s�v��J��� �-��EN}�*��`e�g~�ޣ�Tz^�i&߃k
�;N��޸���O�<cbwOz��i=��$��|�VU�O �*~�=��wǿS,s���{{��/��32HA��$$P2>�g4�� ^ۏ�e�p&?���O����}�nD�2��3B_e��o5�|��X����O=����jg��T'8�t��Kdx���HM���7`�0a��v��7QE;,!�q�هD��dD>T$P�ľD��L�y����m[-��T=6�됿ӛ��_ZQ$9��F�^���NF{a,J��Ą��I.�E5.~�	��&r_��s&{-�4���2|2t=ɖ8��3�Aڌ�9�����@2�5���8��;��_��<�+q?��!)�E�b����藄��=�Y�|���fJؒ.O�@$!X�/�"��vajBT[SUB�<�Ǌ�b�$��2?���Ʌ�U)��X���ܤ-np*Lʒvv���͆��,�!=��S]������.��|�GsVzR�m��3ާq�τ� h�����K[bѩZ�n��f e���!���aB"��Û�x�6R�
��C?��S�]���GW������j�A�$�4֮���jEA��#�F�JW_Q�YyR���9߬�4,D���V�v=M�>�=��|j��ebzZ�+~! �d"pn����ꁷ�Цe���FM�v�/=a�y1QmE��Yxxq漿a`����/|ն�/�) ���%�J����w����:�޽`c� e�r��HV���h�0����4f�_��G���1����0j�{;0%&&�/#���d�x��E�C���S��I}C�����}�#YD�����u��*� V�������i�7�q���-]S���!j�"J�
%��w}P_��<���w|]n��S�q�lB�|y�6�9��$	��7
`Et�!;Z���s:�5;b�Z�:��Q�D�����ӟ���<͓�*a���c��g�������(�h�Li��V�5�w��W��C���$�Vp�C���΄�Z����bc�N��/cj���F%C�	x�|����Y���!n?�)�+w��޸���<���42	l�J�l�AQT��k��0��ܘ�.a ���% �x������M�w�=�#�~ư���k��ڪ|���ƽ[؍qJ���� �O1Lc�T3+�K�u�ؗ:�N]��cD�umC���Xԫ��=C�\A�MD��A�_qЖRD�В�"kv���G���>>��ĩ���%�ޅX���O}�Q� �� 	�i2�n},��:di"�#Vu��dĘ'e���(1����M՜WdGGK��/?�ج�C�19����C2�����m���e	^�n5�>�x�#�$��/��wi�E��0���󋘃��?yl[�dR�[Y%����$����k.ܼ���MC�$0A\;��S�L�t��ưi[)s��M���HWPP�����U�
����KQ@�܂q�� ��l{�}:�k�"��` �����g#�@�ȑ�[]�Sԫu�c�����Œ��>&��}R��'RW)��Y5���b�]�	��C���JV?����"n,��j7��=�\5$1��Dv�&�I^K���M2F��Wv_и]"�	���2SЎ|����Ew�֜���қ�g�$�Ӹ�m�(���s{��R�ECb�/3�x�J�$F���J�����uH�u��|����j���\d��A���Y�r����8Z���J������v-�_��Rh�NPѼͤX�\���ݜm���c)3���c��;���������.ڹ��>揄>�&]٪d���FIuEm|�tL���>j��b�Ng�5��yK޸Z�#f����{���4�(1:�%���8�_����=�5���I;m
��'�P�HڋkZ�v-\�u�!4""a���Uz���:��M��#��~v���J���.6�KKt �C�\�b�H?��Ks#j�(�I�Յ��RNFF����-�Ĝ�Z�q����2�߫ݨ��Wͤ;4�+�������V��~>h7��k�Ң��r�J*6�I���1�Sn��S1�������~+�.Bm��M����S�uJ��׶�N��;����#~�.n�<������~;=��<�x��������n��.��l��c�;���y��HO/Z��UK���/J��oY����i���%�w=���7��cT������{�2�bs��]��E�Έ����@��9]�?z{��@��r����N�OŮ=�9ۂ�>��^'�uB���u^�q������Ԏ+�� �.8�*�$��o�$V���8��ʯ�NO�:�+k�hR�lB�!��~5���=7���w^�
���Qu�×^�;����e`���^`{i��%3l�n���'&�(q�am�A��6k�V$ ��8 %wn;�V�̳�����}|���Z
@�G���u�����ป�_e��x��� ��Z���t��곯�W ^X�|L��P8 0�ǫ�̙8[>_���.��Lj����ȥ�d�@=οa61OH�R��_����r��kbIK�J��;�����/����w�d`o�l"B�[qg~X��Ki.�����0@��o^8<ɫu돗���$>-�g�!LRDjXvϴ+�@	o���FI	�i�y^����xnf>7����t���V�����4z��R:[����D���6X?�!���r�ʢ/�
�ƖB�P�������vY���vP�M���9�������:����h���Q;��|�OO<�sx�dm�	�Ɨ�F�_��t�\�*>��34C�H3�w/ց���o����#�A,�]v�[���#_Y8��-qb���=>��CG�QrJ���м����{���87�w'�+NBxh��2^���l�=E�bO2�'�B�)S��un�(̽e���;��;�*�yZ�}�ϥ#Ę�n��

��O�g��cc;�8��;���Z������|��u�=N�&b��{sZ���6������Iol����Q-E%%
�-f�(�	=��Rz������|���f��=rg'E%F�~/����U��k(�ۑ�����.�&��)���9��<<��W�Y� %��8́��F�<!��%�=z�����F'S�%Jp'��K/�8�KJI��$�0��d?��*���>��S��1���s:�[���A���}��/�w��DE2�*#��Z�2���ʱ��֨�^s���[������Bl�ջ2{�	���%��l�uǂ�%���n:(�tD��������C�w%�N�z��(�ꩩ�jU���`���:p���l�|�=E�~����P�U�\�)9��Y������g0�Q�LNV�q�����W]��J��?'���ݴsS������gf��� ���y��eg�s!��/8�.����꒴6m����������Ӡ<�-�.<�p�	�;����մ6%�ڶ8Rp'm<�X���u^EŨ�$a����a�G�&U�|�C�7�2�/���x�M\�U�����é�4�Rl�On�IX,;q,�zBo,[ք̵�z�?��/��u�҈��������ޠ��^ ����%�ǒ��G���$�|�'�S�l+� �Ó9h~-���sR�?@���,�l�Mx���T2L{��Rc�9�Qy��x]��WV�Uo�H���B���hhi�2*��Z�ir;�!=sGz��RJg�.�O���;�W��l�	����y��=t(>��È�3�»w�&��BB�W����/yoc\��}��r����G��b�������N���S�P�>Z��˧�46N�?i�IR�}�R�`��Fr�6�to",�8\����?��纐=3�k���y}��*$䵗����#�Ǔ'�5�d����8���W��)ݥ���ѼSJ��aGx��Ir,ED;�����I���C��7�X�����W��.Bˮ����b����T/d��rp���t�;U|\_/���� ;A��cc`��GeR.A�ov��d�y�)vH�Fiz׽DK�D����L���i�pi:�q�ϟ?�J���yOV������2�E��T(CP�7�Z���Ozj�������Q�
 ������=M��Sݝ2Yy��]���j,�Ǐ��>�>�w�{��L�^N�nk�F.9B��= ؘ���↘�|ܶ�k��F��u'�k�V�[��f�'�$m\(��`�m<�%t���B�{03�_U&�8.��h�A�� Y�ˀv81�z�<�(���}cƺ�QZ����֤���T�yӳ��J�Td���gxcdw"VXNN��ǟ��b/�?��R{��O�ёǽQ�‍���Q� 	T�T���;(r�c���� ?Y0[.T��%��1�t��e��Hz:��QC�_��ͳ���0�wZZk�I:5���o�T�XYX`�����U���߫�t��%�GMe�Wl9^�|�5���!�����Ru7m2�)�&ks���+�Q�<t�����6�(7d�A��1�����+t�ur��m
��W;�����|�{���� ����_f�wn�}�!��/(@ڨd
�k$��()aifw{X���V� �av��xh�%m���P<����`�B�l���<���>���kk��z[�M�x��{n/8N��\\j�[�p����rb`����R7o���'|]�.X�m�nШ.]�TdMN��Vo���u�O�g>��/����4e/����q�e�_�n�|�o��R����'�Z�K�͚�򌠂�	�p4�����_��,�K ��$H���e�V��k���!����	)LԾ�U?i�hC��MU�y�
4�bׅ qppTl�L��S��.��#���Q
�_Y_+t54x�+����������5h�PHa�9�9i�󺻀��`Q6��ဖ@",���_ c7j!uss�zt��h��@"bϚ��Ӏ�N�����v�$|����O��vs2����̚�fC6C�:��\x<���s���|p�ͤ��F\LDfu2���"��P�]zHW2X�(��_I6Aw���p��ap�
�v4�|MO\'u�]H��~q6)�Ŋ!ٺ�9N}�B���O���"_)�A�n�B�.�肵}715�ݽ�h&��F��,�<���� ��9Jlr��|h�I �;n��Ov��?5�d��'� ~�DAE��M�$� '������E����� q���"H�T��c����͗o^�*��Pq��[�Io7���Up6'%���')l8'�fWSCEC6񾰰��P\�4������x���yCw𥚎}(�3��1�.�����m��I��cq�	�g��D�H�o�om�3��e��#�T���M��*��B�N4��ݯb%.��[�^WU�AH� 6C���`gi��	�s�ϝm�U�c[�A�6! L;����1��+~tC�:�J�����*Pd�? �Ԅ�>ָ���1{˯��0� +�O������B+�Tw�����\YN�髁�g����C������,������:aH��!/,.j��y���b�����I/zȌ�'�۱7M�b����%5Eǹ�ǹy��Ff�[$��>'��DҒM�o��(>��o�/��Z+I�\>K�/�O)��+ȱ�$��W{ �e�\nm8ɿ���E���T(���w��,^ ����h�I�Hgam-!Q��3���e���-,?�~g�{ f`� �Ė���o�?��Z��P��~�Ȑ��aS���bHB#F�N�^�Ȱ�L�E�.����M3LA���`��L {t�"�[B��{�(�n� 
��a�"����]H/�p5\��'�mE�L�uS0��h��`�u�BT��Ŵiٲ�r���Th�1�d�c#�pk:#�&H � E\��\�(�N>0f��?� .o�كOlVÝ;}�5"_m�q���B�ؙ�~��T�a����K�z1S�������Y���y��-�l�֋>���?8��gB�n�D+�cɀ��6iИB<J���[�w*�&dX(���z�g��U��'-��>�f2�.���"������.|����0�0k`�N�	h���ð�������MOO��٢aF�6
���ű��6E��1z|�����?M�络ɀ��O[\f�`�:ۆh9�x�Q�`�g��2�!��}N�4�F:
�:��z_ZzW�콼�yh�ye������n�Y��} +x���T �.ŶhhkG�Đt�^� ���t0->�\{�D�x%��6�@-T>���ewP�����'c�?��//I2���pt*�:���3�K2��(�{pၐY��QI$�X�{��^Ө�}^�t����211�+Ӯ�7�ɝJ>x�����J�G~����C���{A$N�жz^���`gT�cW�����χ�'��(_� �*2r���,��� d�M~��_�<W�Zuf�!kG��zR��uz��5�x�&�O�p����u��ʊ�>)2T���+~��7�� �;�1�z�2Y,(��3��4-Ez�2;!��Ͼކ`�|�Y���C�v���og9��y�s�,uaf ��;�͘c�q�\�Ď��ǂ�$��H�M�Ae�Zq�s��z�꾧���p�U��SV:$@U�쪾��[��Z��ӧ�OC��L_7r������d�����|-��?��{ÿ[�KC||p9����Z#�o�\��	w��:�XV�<�O �f:�j���&�<��L�,�
n����6��K�
+�-Bm�8lϜy���nֈ�.I@NC��;F��W_�a�E_�����dN�Wqr�8��Zq��wvb���֓L�A�mVz��C�H�������#~P�ٽS��;�cY�%��v����T*��$�מ���t��O�Io9�0��{[L�����)Pʐ�q}��������T.���M�i�k������	,����48
�$7��F��&}?��g�`�$Ӈ�N(�3���F?{#	m�&�G�Q�/��w�o�~���
��Q��Er;���1�M�$iiY*K`cm-el�d�Z`�dfG&���uG�2d�,���&�P�ĸ�_��N�Y��A\��`�̘�l����x�z5z.WDDĴI����Q�h(!iPjm�_����@l,HQx��6ĩ�g) ��W@I+)nr��Nj=?=&O�����嗕͘��H��13��0N�B��Us�K0pE�����oya *� ��#�E��N�g������M��e��{&0�H 2���i�N���S�U�fl��^��;aA����ѽZ�DzY�H&��[��h�Íd
�'� .
�R���ihh�P���p|ײ��vj���=Tl �����^�_�͖
�l��wA�>PQg�2l)�rɟv�u8���O+�އ5s�h�:�D\�2,�VE�ۭ���0�V�PN�ل����X��8�&g���iK������uu%7C����XE;Jr��?{�f}յr]=&�z�
�� /0�����W}�L6��� ��q�6~	�А�[|�P�����Jtm���Y��Z|����`�:��.WU�y����V���0�Z%��Ԩ#�\�C#7�������� �v�rc�`�{>56�ӽ��O҆5_�������塚~�|)�����vL?�^��(ϟ��>�Z�I��ٳ�IU|��I,9��%B ֊ҍ�j�ćJ���o�oNM��p"4޾5ӣ9Y�Vaē��gχ9���b��OL��k[�]�uL���n-!L��'S���HK��5�=��=�# q:yT�h4rA������r'��΍��U��l���"�8���!�����9��qN�8�kh?�+���g��K�nԔ,�O���HO_m�~D�����͛-�N��_PP�?^����d3v��y{(���}q̒���ɠ�����c&��z�4$<4�����|L�󔶷��1����2c�[��E����������t��?�қ�n޴,6�G�V-�	�P�0��q�;kI�;����~�f�`���$�Q��\��߹d^��k��K�Q�pU�kkk�\:� ��A��&	1��x�`���&���O����W�Ũq�mMf�֟b�1�(��k��z0�B|���#p�6.�_�=:�i񺠔��G�������A�6⹸����X��6>K��Z�U�K��0�֊�Qgz�&6J�lU���S�L�v\,����dIX�}��=�`������t.�YǙ�� �m
��v�F^[��<�X��Ko�]8�P�Ї�1�1T2M��o|O��1�o�=�BP'j]+��y�`7�T(��T��7qtTT`���rB��^�e�[����P:Z��ckN�_$���.7v�?�^�K��� # �*�:�㕝*����n��N)�܊���֙��I@�6/��^D�:�u��4j%g``�lz�m���!|. ���;���2PV�^�^�C
���!���>�LZOa�A�;p {����ūsJ��� �#>\�Z���PEN���u�<��×�^=�5�g�	*_�M{��^�P��C �0�?�>�Gkyɹ�fM/.Ƭ���'B����2���8����c��3�wGxd��4c>���N)��߼��� ".&����,̩��F��J��<L�"s|��f���l��N���r�_�{{{{��:5[A6p23ix�e���eq�p��w���+�,�Ep'\������A{Δ���:tt�Q�H�� �:~%�Ҏ�!��@�Ѻ��	�?'��_b��IT�N��~J�l��y.����r�B� V�2����" >�ޗ W�t*+�W����z��xC3���R��k�ߚ��A��zl(�R�l��&?�:�!�=Ի�J�'|@ť���nە�'(o)���O�K'"^[�o+'��X�65�}-~�(��@��u��/�텽��L)�O�=��8Oy�ǉ�O���I5ޖ�osLĞ���ݔ���]	@�x!N��b������Yv���"=%��f��E��jI;O@��K#���8�e�;x�p�K��ï
���+q:Yt8�@P�Г!\C��k�R� ���K����p������UW�����ٙ���f�I�uG�11(�(l�0�zyy9C����]�ϟ?zN�@S?�����>ۊ~>	����RB-O���29�����xo���akz�������F��Pk�_ �4��3�f	�qǬG�J����h��1HI�0E�4�X�L.�f�p2�G��&%'�JQ���y���=�U�jط����x]Cø���əX[��	�Ҙ��qt+!A�y��)�Dɪ�1���s�;�_~��N|EJ|^
P����j3i������Y|pLp)�g@|��~
�-�<��>*���)96�Pu8Y8�u�l��A4�׺Uh�Ʋ�g
��D�r���Դ hǭ.UqO�N�?L�;��RC������)��j�Ԑ�Ⱦ���>
"9���d�<�h<�ܱ�p7�*B�jI&�Io@�;�%�:\��$)"a�'&~�fec�6��I��y >��[���p��������H�����?�������F+�;K�	1��M?����c�: �*��?s�s $))M�0_oG�y���ǏZlcTʪ�5�(�5�Z��!�~�#eg`>bW�>Cx���/ڧ��8+˽=��g>T@tgt�h�~+(@�uT����gn�t
	�r~~b��>�u�޽�k���g!���(��^>�Y(��8��t&�<��2�D3B��jI"��W�o�u�����m�f�"��
|<::Zv϶x���j_]�I7M1%�#���ę���DY���ޢ�Y�=R�������������}�+�V=�{%I��=��������J��ᣝ��8���	���t�_�hղh�BX�fpW�[���Gm�I�3ƒ�mr��Y�U��XW����W�� ����N)׬o}��f���X�~����H�K����B�h��0$��R�W��Ot�G[�b��g���؏t�9غ��PX#2���ٗ��\�&�k�J???W�Q�4�����I%�}z���ǒ����v!�Td&���(�F!Z����..|����֑���O���X(I�/i������+�SJ��r�]�?U�wr"a'6�WN��&�H���~��	���\{"���?�����_�:�Y���Җ.����h��a{�ژ��� �y�����옓���mo�䫫)� B��խ�T�όe�>�c�a��vd������ �q��נ!��엫���8�p9DҶ�=f]�6�['8��3D�*��^��=p�/�0�to�㋥|�b%��H���pQGe)P�~���= U�dC ���<񰱱!�[���0ѵ��1��7������-��;2֠�a�ЋɆ�� >��~�A��[���T��jHv��(�c�)�&��KA)�����k$~(�����>lm��6�[����p2Ӂ?������HM.�߿���Cp>�R?�� 7�[��P˚�#��>�]�X���	Ϸ�#��/x����.ӊz�����B�߽:WA�q�aPǮ�q�bwsy<ୂvZq0F~f���'5�����c�B�����I4��?�3'JG̺�[Q�A��a	��)伥n6}ju�V��"��$�kě8S�v�0�vkk�d��?V<���M [NB�Ԋ����͉��;6�v����ǍC����71"�So�ѻw�6^��:��3�I���-�@��K��H����txq�N�sՓ3�p?������r��\/o�
`@icgg7��O���V0F���@� �P4[^_?�t�77���� �4)�����Ծ�ǽ@G{���SS��'�v^��G���.t����B�[�^�@_��|��Y����`���/F�O�Cx3�欢UG�ĥe͞��̴��WaLƢapXX�X$��Q�XNت����)&��eE�é����9���M=T���΍��Iy��`��	A���k��f�i�op�&�Jo��	��F�(qܞ�l��D�8���j�C]:Y)���f8_��L�1;+�/�0vw#�d�����Q�B��ߒ�j�t�$�����tZ�n����{{�/���ǀv"""؍i���7��͑Hp�?.��PJB�j9.`�h;��0%�7* 1GJ�J��Xsb��NƉ�����_wL���1��c�|'_&BU_���,�X֤�FMk�/"/��kt�teD񊚷\��_r�\3� )_��Y�[P0\��5�����rOc�M@�2�� �+���ߖ7G����-�_b����m6�͇��,u�(�ǂV/�����UK��
xA�ݾ3�S��7/	�̬��3zB�,��7���17� ��%��h�iu����ܼ.�:�q�{mB�~/1�@
T���HZ;�E��lt*�<����ĹOJeҴ�\�
�h�!+����=E�����Y���Y��q�sų�&����}�g	ކ܎"vz���3����jfD���5�"ʺ/B����%����d�n:���NL���:
���7����+-���-*hNB�Cpm���
^ 2F~�~����Z�������M$���q�@_'K�H�(��0b�'�Ѿ��|�΢f~rf���z��K��4[�I{���ݓ�co���\�i��!�7mkT[0��@.Ƣ�3eY�N���h)���2�n�,�ǝV�w]�b���0�	�4��`�	Q�����efv6���@l�x��C�U�Eյۡ;�Q���NAZ:E@�a@@JJ:�i)�n�����S������w/?��̙a~{=ϳ����g�U4/�t��e����6X����Ѫ"_�E�KJ�Iu�t�oP�i,�K�Ͳ��#�بʨю��^���t35d��|%~F��[��Ǖ�e���Ҏ?�B\hx3�MdoO<�!ea��)otv�u��ʧ�#;M�l;�,�K����˦�r9%���p+E6� ��1	\9+�Ayt55���o߾���_;�����T�S�9,�4��]fB.���@��Lkn���Xy ��}$�gy"�L�4�pO�of����˹�y!���Bo1��'�����JJ|��!T����#����"�o�*U��l���$�e�G���Y���,�qRĐhB���W��9{�9�@����Ê���.YG�╈],5��;;;��bәb)���?~�E��>4���,����2�ߧ��>�ub��B� ��
cXD�%�E�9�%�3��3L~<c,�	�ktʖ�(��拯��&Ya�A�vO����BV.��H7j+��[�Aʼ��O�[�,��U��ͳXmW����sk���k<����'ξ:��3O`@�`�B֛	��M<����̵H.$�"�^�*���B����rXTʹ�V-���`2&<{�/���l)#�)C��k*�_{َ�g��P �mh�N�&t�S�>��mP��@�����D`hd�82&cd4�s�}���Wx�7�䐐ɦ���i�O<�BN�����
����}i�3]��O��w�NP�W��K[�E` �'�m�M�ˍ�0�}Q{�$(	����S��)O ��Y͸A����$6˧�t�z������@�yv:�$�k�f�&�&I�j���:/����������dz7{J�����������~�i���Eq�E�\�pQ�6�ĺ ���p}��ל���û����V-d��IBA�h��Y��wc�}��؃�V����$OV5�-�2�%m$hW��C�zTQ��1�/�Pl㮛A��G����m�o�	^��^�x]���&�;"�P����X5�8�wO�!� �;CCC��rk�k��TL��r��9���].�-:�j����Z/7��R$)�@���g��U��̳|n�g1��פ����s�,�|r"��wx���*�O-�*��:�c�=[gOΐ�xUPYISm�����>���/tG��U��y�,~�0W�G|�/��*�2D&7>L�c:��lw��iQԲ&+`�\K��]y�ryE��7鯬�YW��WEAc(!ad�(�y�)f��+��`��e�Y�E��P���w���Qըh��E?Ǥ�šwR�8�>��j�E��C����X���Ag�&9�Uߟ+jC�I��z���mQ�V�I}5b��9��v{�����m�����(�go�6n���G�ńk���6���r�Ƴ|��UO��bs�Ȝw�?�/��G)4��
�b,K���o�4q	������J;5Ʀ*�����@��nft$C$i�4|w���29>Nf������5G�a����v����˩�����S5�l>��a%Vr�7��W��dr��[l6��փ5k��J$Ux˚V����߻��H���k�mʂ:8�1x��V@�N��%9�?4C~7K>��f�GV��E�PG���A5$��U~HD�����rE�FUh̛mf!Qy!"�x��IϘ���Cj�Kxr�io�!IY�ɐ��F��D�G����7��<��|m̊3�&�Ѵ1j�b|&*2фpey9���5��K^��E���h�(d��9���р���º�T����c�<�o��$�(Vy�ǘ�++y�nM�^�k��pKR*�[>Y�����Qؙ��>Bx��3�M^�J�=�+��݌�둌�z�����E��R!q��Ҍ[H��i�y����z/� �B)Nc^ � 2@�a��1��=A�(��٬,n�}<�{�����j²d&&&նUm���$����W�3�:J��c!�V��,�6�EI6㻟��X�|�J�a��::� E������6 �:2j���QF�Z����~O�?�5�3�p�mC���]�T�ݔ��Ί���gqJ�����a�އ���_��������C����k��n���P���_�KE�Ҷ6	�G�Fq��3��U&�]h���X7�5�_�ݲ�)���[9��� I�L��d��
p^Y�����!eb�I���"_Q�����,�΁#��w� Lyk�n[Lݬ[y�7F�|�|3�[��P@qL��/������&=[��_?��l`��I2E��'ě*�e�@g��;��m��m���2�K���J����!Q �����kFYN2_n�(Od}��5V�����%�Tп*��^dUc��ȭ���?LR��;�'t�����>U����NV1s�b^�9��v���������Gd0�����j��"ҙ��#z�ȇc]u��s꧗X(1�$$Zlv^�zT��:Hf����~�n�q�Ph����?Un��E�IT��m~�SG�����R����W�n��wC�K��R�q����q֓�� ���Ӕ�k*�b����������A�����qׯ������U���V���v���-)���C�v��m��>��tG2��"F�{��Rbg��:��gL�[���r ](����[�uo������Sb��/�8��r2mlKqÀ�1YT/��^�pzydTT���Wiuӳrx��P��2���>�x�nM1w�b[^Q1z�G���U�~$!'�����9�ALY_{������[�*�fKT��q���M�o�&��n��bw��{�nڲPI�|�n1��3�[�u�.���o�_ܴ2?f�d~*���[t� �D��>M/1@���B	���A>��`���*���}�A!�1��x�|5dgs�Dp@�,��������,��;�}a*'{gg3F(n���9Q�z�B�Q;|��艐�Z�e��-Y��*�T�A+P����m��Q������5����߿⦶ō.c�qc� Ѫ����}#�<*�>[���0lu�4�����٪_��./�����)Oi�ٯ���6[ﱗ�i���hDm�	m*��K�%�,�d��3�,�=��o��m�}�L�D �T�;�*�1�oa��U�����^�hZ)�� ��9�@�����-s��o��2_#q��y�1�����$�4y����{�b��0��Z�7n�x��4���<kr�v���xG�b7���"�B�/�L@>+���#���GN<�D�*Z�)�W�h��?j�8�c�233)�N��F�$�	xZ�AM3}PaH����>�b�����&I��s^);�����.輄�=�U0��y�,�ɪ� o�立��a)�Ksˌג#+uDŗC����� 6�?DZ�m�29%%��^�}�7��^�^e���t�۪YNQʒzz,����U�d�vYC.��RA6����b���  l]�	`��APdh��]�K k'����������i�y����@�sTw��%s���Y�*Ǯ�����I���f����]'@��j���߱u�M���*<��X� �!á�J���Z��HL��Ynt�(�#v
������H�f�LNM]��;�^\��{J�X����w
���}���{���cғ>wt ��Ϗ���=-����1,Z������������7�j_Mܐ?��/<��SZ��,����I��=
����7Ui�@�X��`�U9'_ �{�=yYyH�CU�8$A��76��N��4�9A}�Q�"�q���s 9̙�;�%�OwP��xz���o��]�N���Wa���A<�q����-")s�����v��g��KxO�@�V��f�B�.���Q�s#��:9���.����\�S�Aƨr����g%�������4ȵ%"����7���"3�?j����-�M���wY���y�?�IA�ʕ���苾ڇ��wkg��{+�{��I���~xs�^���~�)�e�;U;;8��:;:�V[�>z��t�<�����+������,�Xm�)GTא�����ӌ׋�qQ|��`fy!�<KA�{���@ӱ�4��"`�7\T�.$�z�T��o��|��SQ1�2�f�N����iR�_�ψ�-��͋>���H�����~0vU�QHD����-,�h� �&�<�+r�V��c.���Px�O)?}�i��*d �qk��-�p�a�V	("s�{J��'�x���kB<�:��@�5t���5��f�����<�?M��\�D!�v|��� ��a�sވ�\�/�ݑ���S4"q�P	)�j�S�N4r��0�����>bu1����~	���GA?� �sD�W}��<~���TA��z��x~�aE������� ��W���mm�$*���/��S��ކ��
 �錏��`4<�&pf�[[;�����ގ9'~�z����pm0n���W�LQ������"�61�W)/k��Բ��:��9`1,��t�D{�U*MRP�C!�k2ﲛ+��N̩q~rV���q��%�(Ѵ�d��=wtw�jrA�c�Ru��) *u�pwFS_�9avt�>��dn�?k%�������]���y�XM_m��Տ&����ϳ�WL�e:3�Y��S�ٖ���A�,t���[D��s���Kq�"���Sn�5rG��9w�ƒ��-%����K(9.Q#�O�.��D罭W��6ӕ؃L���hUV��o�n�X��$3B[�]*��=�Bܪ+mYZ�_�6�b<c�ŁRAQѪ���9��M�"����@w�v�Y&p24Z��M����!���;�bG�Ż
N��W��o��e�b�������3�MM��
3O�G�%i�K������.����z}f�r�U��0Ta_ ��U��ؓf-�Gl�c�'����l\��68���?���%v3V�l(%a�ڂyc{\NE�Ԓ��^�lp�	�Yw��f�Y���ً�l�e ����Wr60�F�i��I��M������Io�K��v`������M�`v���̇���>����_��f$;�p�T�P�1�\���jlg0q�6k��X���&�9���$X��G���Q�KEl~+0�]6�)b���j 7����hKJK���?j��z��RY�*��az�8cpgzH��޶�����Ȅ�آ���Q��*̎���I����AL	{���+>�z�}���r|���ޯ�	#7a����WĿi� ��DuD�!`�j}�B�RQ�?.U�d�@����LlΓi>��⚡�Ƃ�������y7��'�*�F� ���o��%q��? Y�o�����&5N�^]YY�z���+�:$#���,�ϸ��h����د�zߩ�M�2
�v?��+��i˼���F=	
�_}2�g�y�d�������i{�g���\���D�����;�Vػ��k�%e���on4��\)���m����Z������h��6��P)k=M� ��������Dc~QQl��"tK�̯�x���rE��>NW&oФ��2�A�Z&s"�VG�w0� ��� 8pR�AwP՞(&�ӿ��_ۤ@ÁmY��N��2::����s����5L���\u����2��QS?9��˽·S���v{?��[nv��Xgy��A��=��`d,��}$5t���jc���tt3�c���Te(p��)O+He�X�B̗�]���d0�o���a���B`1p���[&��
��V���a��R��k/UU�Z��ᤌ;�X{��e8{�1��{���DE~4�VMM�$������TyM9j�=n��ݥ�ߢX�}��\��_R�sh�ْ= 3�
���9f	��;(��Zm+q�a�m7r��ˮEp�X^\�7y�Do��5��Kuˇ���^B66�Q'��xo�}�#�͟^Cj�!��=����J?�E�o���]ۀ�#���F�I�&a��\$ع�i%��WC3������RI�5]H�e�`Q����z����kb�K=/}}y6xw�h���WSl½�,�����I��lllA���E�(>����yZ�Q~jj�1�w���,H5��f=tuj�{�v7k��h�&TH�l��'����:<×��?���y�ȯ��;�*��Y-)!
�������ТD�a�n���(0$$)�W[�T�>���=��̹�8/M=�e��8�uK�P"N{ �74~�_E2�^��l�>��!4j��|ĲR��B��z[�&��2ss�*a�K������ � ��Ms>��qok˶�E%���U�#����w�]�%��OγWVo��Rw��$�?s;�U��!���sk�����yVE*�I�����..��?
u��0U��o����2��,�����& ���uR��&ft��ԭ�����:D�	�6"d_f!Ý���ܼ�}ie2<�QgV)=���3�)$m�����G�:���&��R��C�[o|�ī�y#�SPrbp�C�����	O�R�CܺKtJ���3�3��5�����U[�4�Gؖ��(�$.h#.Ƌ̖&v�5���s:�$L�≊�N�?{�D��͹/��qy��E�����ތH'��6Ӕ�%����8�	-T����$|�Dܺ��,�����,��" e����SeU���Ln�uә���O��imjV�Ԟ8���v&{�s��x����%��;�J����L�3�����P�x�~��/C���B�&�};����C�N��US�#~���@���S����ߪ�n>�suR�gV��W��a�9E����i�i� �ҪO_噿Y�x]
�7��g �x�u]a���}�z���egwMZZ׎�"��ԏjT��s�s\�>�++t�FFV��c2��;�Z�^:����8c*�,p��S�6h��PZф�V8+q��u�j��D�i���R1��� ;v�%�c�j�����Ԧ�ȯ�T�+��.��!��[�e��ᮽ�W���An^�:����<�-fv��\�	ڗ?1�{zx8 �<�tF�w�U*V�W���h������w��X�"$��s��vٝ+n���g��jy�ʕD��FY�ZQ՞�!kt���w(6azhh�e%��
NZ�=��|AQcͣs������hF0wɐ�#	�A
�q�"�W��@Lp��*%�J��0))il֗�:��T�GjOOS��YI���y��#t��H��I�49��Oߡ{���5X�8C)��f���GR�L�w0q�E�����h���\4q�������`jj$-�/r�rT&S���u��5��A���a��x��4q�ɠ���hn��G��;�|	���7����aJ�s�����'�ݷ�@�6E�S1s�Xbm��/Y����7::��$��������,j0֜�yxP^^��n"�v@�(��wݣ$1$F�V�u�_痮6Sl��_b-n�����!/^J����0Qd�PY��_��]|�]���b
�W5�A��'I�wy��R��J�s��O7U�pcJ��q>�ӿn�B�f�I6���Q�5���\K���%�Q��Q�]��|��F�F�� ��yQ5�Mc �o��gb�����'��qk�ed�sENUY pxZ�a$���G>Q`��}ծZ�"�Ч� Xߥ��P5���q�'�p\@�k���)N���w��Q:=tx��ʶ�w�W._�Xyx��
�C�^�A�HUg?�s�$��"�Ξi�nb��KQ�]�d��"r�-��]�(9!��?'���4%q~oNĚ? ��j+��^\6Ɓ $�"S�5,b�o�r	d��i�x�H&�0��t���0�b��2Gȅ�C��%�7H��`F��6��|���}�ԟHN���ST����L9G`��G�p3X)����j�h�f��n_-((�-���0�?}�e�"�����_��x���W��ͦ蝍��n���lBi�{��qZ�݊gk���i���%��������.���33~z��6y�b�EH����=i(���c~	���t� ��i�%	�Bf��b�[�|�:���݇��t��&7���XT��[��\���(��B�ce]���J+ ƪ�N����S��2�^4�q/�޳���ظ�z���Y�a;Z��'oY�f���퉉��_���~��N��Dǖ�+��g�Ǚ���P��<R{�&v,����C�%KR�l��K�Y�a��tВei�T�����[�����wR&����!J�l+����
X��Q�*�����s�S�c����#`yy�Oi`L���R�
M����V�h�H��Ev�̢�X��!�����m��s��VkuF��	�=c|�-bu4�>�*4y�&QM��DH�>+R[����^KL"^@�Ҏ�_&���U:��G=���]�
�h"����}�O��,��q���~O��Y?4#�9�2L�f?�E���S}�T�	�é~���-���p�1�]����7�"OY�2�᮳ �dZ-
��U�� )4r�ve��!�Ѱ�?	&*/t���8�e�Z<���<�A굱�fNժ�����c��,�|���N�Y>*�-�G&Ӫ�U�y�E��W$g��0& nq�E<��e�ϐط׃�D^�K�T��k=������Y���@�r�A*�^��� �����EJ��;�Å�͊���e��}�_:!�w%�]�gr��.�l
����~T 
�����ی�H��V������'D�ǒ8�V2��!�Y��F0��bm�9��1d���Ox��3-���t�x�U�W](��>H{��*��,}�"C*S�;���.�{y�aܜ����k/H*�|���r��@�KW�9IZ�HV>�"Ǿ������TA���c�#{ۚ�A)�Y��߾Yg�B���uwU;d��M�c��[�h�*�t;�;�M�`�p���S� Y_�!pJ�@��������=*�z���;�� ����q?��nH6U�Gxnn�2�ά���
K�.,��[�T�h�z\�P̻�7��E��k
����s�H��ي1���Z�&%6~��G����x;���[��r�fw��c�ج!!tu91f��JO9��H_?�Z�-Y��|/��[��F,��1]��F.��	���P���!@���I�����n�����ÿ�b����>_���8Yɱ���u�e�]t�l�����f��9Ӳ�"�����P���p�cr����|��Qq�5r�l��{�ƞ���!��+�`�b��6���a	<ß���mf0��r�<�����Ra�t�H�8N����aF(s� }J%�Ye�����60(ׁf������cУJ\��PH��̋$��T妚����k�A�t|.��Q�h���ꕀ��pl��FO���U�f���3�4�����	0�Ҥ �>�B��$9MOG��ϟ��ҧL	Or�9��le���Y�#����3I>9�՚8�	;�����R��3G�u��Z����s��m��aɑ�	F���T���Z o�W���n��}V� ߹o#�J\�j"mk��6�%G���bG�w��J�EFXb��͛v�[@�cng߰ͲE�k	��[v�>��g�}'>�����n�O;vv�|5Q���a�$��Ɠ���RQc4�j�蒱8V��ҀQ�bj�$����4F��5ɹ���Ꞻ�)���/??#���ӧ8N�m1������~.m+��{'�O��8�a�u���M1�N����BSR�=�}�Z~G��-�nӒǓՌ3�;���tP����:��8i��#��uu�,�5�f�3r�Y �Eb7;������B�!�}��N谏Mx6�p�(-$���z�If�G��|�44D�I�@�82�px��m1$�H�Ơ׊�U��3tJ���A�Q�xbW����S6U��8ΎvZ'���o2�������L썋pth(ڬ�@7rd�Px��X����y�J�{�~���3S�:��Z���F[��O59<�;�5���?g[t��o��$S[�r��3#�9��t�>>>��W��zb��J^Sβ0�f�I�$�6�i�:���o�~�Jb��A��~!mg_ ��a�^%M�QuM��F�l	��9��R�.^�V��q+�^��:1�Y����`�z3&.�Mf��Ɨ�����^^���h��R�kܗ�gR,$������P�iƊZuՂ���`��!�
�.���z� �� ���{k�s���^���iD�k�\n�#�������h����{��
�> h���!�<��U4s����2����A7���9�}>_���
x����%����eޓ�:�v/��^D�a.�VUU���O}�0����_�Z��l��U��󋋘��?V��Fv��T��{?N�Z�`�L�<��FO�46O��·�PaT��io�=>>��T$ ������h��\?/Y;�k{q��F>��1��9=��P�eӟ�\B�cY��l�T�h=�]�L�6��ԇ����/W:�8��҇|z�\`���j����yVm��mN�G��Y�ܳ��# (=gEzK��z��z����M��9zV\�>�D�
3 ���N�%���%ϦS�Ģ�'���B�ES�8�ܬz���uu:0���G��������>��I,�/���ާ�'Q��U �jaa�J?�Eݞe2�O0ߡ	�ڗY��Ɵ�,��c�(��#%�xA���+2ss���`�&�c��P�h�(^��6$������������^)>���_���oJ�P��U�a��ˡu,��VԪ�Ǫ+l��9�V��BM��--�0ahh�r�&�o�g;ɋ;�H�~b��ΐH�~*�7/�]zf���gIp
e}����@�L�|���.�)\|�#W�o1>I ��,T��]\Dұ���0����C���v��/y���vUǴ�l�j�~��L��"ɒg�7�0���ec�;�v�+�2��F+F��G�o�m4�]� ���7�����|8ݠll�hى\%&�%�f{�+E��7��Q�N�����dݷ�z�R���2�-�A�
�T�S�(�ϟ��7u�EmY$��]>_Q�t�%Q_q%+/�⮛lu���ڀ0��%�mpe8�C�����k�E�3U޴�|������m����D��A�Pi����Q�'�������ۤj�\�����<�����
"��$̄n�(�fZ�q��2�6�S��L·�.��5`���BjZ���k �jl���o'|4`$y�� NOV��7%1��!�O��~c3℞a.� �
��)�Sⴽ���M��ܷVa�����;kt̘�p����7~����)�/�k���QK��S|%nh��dEr�����ڝ�@���cI2슸���`�FW���k�ܙ�W�>�5�w�x�9�����!�h�s�=�A��~�1w���&��)2r���~��E�=	�(y����uɐ�%*�ʊ|�XI��,�ǧ��=D˯<|�tA�������;ۼPלge�Y�ֶ��P�_�d�}��G����Rµ����[V(�&{r��U5Eؓ��o�8�.f�=,ə�}f�����	�^������i�U�+���A}"_��ns�
K鷬���N9�dQ���層�����wF�����a����U��15�<�mX��l_#t�6�{ϰg�Q!T�e�N[婶K;b�'##����٩�CT0������KnV�{B޼�L�ѐ:��r �ֿ������ݰ��H%�@���8�d�fZ�
P��+Ziܗt�� ��1Y��LG��� ��whoԕs�-}b��%��TN"W�j?nH�	�]��i�SE��~�H��ϥ�����fO�!9��q��x�0�ŗ�+�������>�U������H�ܡ5����cP
��q���lw������2ӆ�B1t�򦥥�m�������S�H)B�p����/0�}�W��	K�&̆;p����& ��a�����}��x-�����
�6��3�^
B��ė���ո0���� ���F�?���@����_iQ�M9]���T＜Bݭ�V(=�˖���4|j�-t���VS��p8��w�a߃��g�M #z^L=���aq,��l+���dw���;m;T����,������;.����a��ϑt{�fA5]_,��n�a�V=�*=�C� ��k�Z	H��Fԓ�(�~��LB߳��\N���
ߪ�~�]�|~�z������W�=Πߑ��e�]�M�~���S;[�����r����$P~�@��f#�*�s:�r0p���Dţ�3�����ʄ*�^��'[�D��N�=�WX�1_�,�y��v42�b���Ț'�Jv��7��8��/���jEV��qO����xL2.444��u������i�M�������Ɏ$��iXt�_�b�H��D..�k#�"p��&�@�F���ݼ���pM��K�����@���c�O��ԧ;�I&8����d
051��P��(�^�Lg˧_�d���1��2�yR�D2B�^'O]�ŗ�/E���GA\{�]g�>~�Yq�Y���f�|�u%���K?�tO��Ǝ������M��~������]Yht����j�v�o�ib3��!I9Py���5��W3��� J�,�:�S�E�U�,�n\K1�ӭ���=���X� m�:}�Iv�W)�]���#�@�E����ox�&����F33��&''u��K�I�+��t\�e47"Ky�˓+Y���j^EB�S���5ٓ���9@lW](��<������%j����Z���q߳���u��Ũ�ҰS�3ޏA�-����;�!��5�k�q%ǟ%���O&z.M"�.}���'�
$Z �A
��1z.��{�Ά� ��*�,Z�@� ��@G�ߧ��aYD�73�͓�)�����˝�.Yww~��nZۨ'_�[�
�j�62YL��CV�%��
��FG���źo����1�--}
�e���!O����r��E��eG���}4�z��b��zgډ_�ɑ�'��T�2H��{^|||��ٓ#_F�R��]p���/�X���#�x�x@�~卮�&3!�Ͷf!)}O{b�Wm7(✇��SR2;�<P���J|Еb�Tr�/� C�QOՇb�N�w�!�<�?� �h��^�^�ġ�sMmcK����(yh�E~��X��*3����b+̉��	�k?��P����N��P��'�'I={F���0��8��!�%F��3�跀�'�w��tٓى,D[\��[�~�ߐ��O)��*�!�h�b9>��sK��V�������y��`�y���k���8������Q�<%�)Wo[N��k�z�����=�[,�В�,,���'��,�\�m>�kO��]WHP0L�������Ϟ;��R�|����&֜?��BE[�,|��PVT�z-fx������p4d��IJ-~�#BӼ�q�n��M��i@�U�]��9����ؐ�����k������sS��������h��m�cc?��j�#����@z��j_Dސ��I�Ƅ�K��	�%Be�\�7} �,4�"FY�X[ki�ag����Xx��-]ʻ[pr/z����94����Ԛ�s�/��L��&3_����T�5_wc�n K�p�N�n���`!7��m��|������mɝp�s�����ߕĔ� I[�89�$R��
1M��ם�gR	��`�a���9ŭ)�j���|��weɋ8�-v�3_���z3��X��NNj@Bۦ���*��`��k�����
��:!E��?�@��\y��v��-�	X�-�/^O�ۿS+��=w����:*4���^&�h�St*'���ziAO��2Se����B�U!'�^g�W<+�%�.�]1��<̃}Y��#/�m0�@�U
�ȭ��q�C�2�w-0#į�ڟw���H�,�k��*�nn�n��U�n�Yf V�'P���'���AA�ԩ܂4���/p
{��\۳�����m�+ZaGd����b����F�-��"����j�'L!R�/���m��g���;ԟ��mj�O^���\b)���ﯢossCx	'O@�d%�jpߊ�,�7��5)�_{�ް�}BGw���B�(�>����{����{@E������0p���]p0v��m��s�
=���e����H ���<&�g�d0�|��%��|d���e1���ON2+���o���l��g�8ȣvŚu�17�tll|Vjq���TUUA�X��#����D}Y�`�t+K�g2�s߿�t=�2��`�������)����:b�	LT�M7D-�}��@�������AR�u��KNn��4��?�%�+��/�y"�P�Bg\�v(�7C,zЙn�dD?{�]W�R��,�PU@H�N(�cE榮 Ӊǧ��`��9-һ���2Ymk^q1Ve�Y��q�D6����rA%ٌ�Q�Pש�����,��B��5��9���^���L.��G��B���d&_����C��J�xye���S�=?����9���|N(�ǘ4��J_͋���X��j��}����w �N�����d�JFFֆ�\k�������!S�I݈���C8�76��ԣYP��`�K���:���q��#V�w��k??c���)O�LZ�ﯩ���ۗ�j�����*\�����"�e�:���a��M��|a��a��t�����2�J�v�>������Q�錰�$^�'�=@L�UV �6�Q|J
٤�0U����bS����^k��ͷ&>��P�������aIN�L934�o>�®/�:3�ɀ���J��y���+�n�hI���Y�2X�����\=��RoZ�i��"=vʫ>���g�GD3��o=:��T�|ܳ_F�q��ez5��Y�@�O�G�����B=�[���X��1��q���]�,#҅"�р�ג��6�F*���ŭYߦ���	
�@$�Q��lؓ�#�ϟ�||�X�?~KG��,\`�j^�2����>��e�c���f�P(�;�E��(�}M��h��¥o�Յ�jY�Y`*��i�<�����A��A��Xv.R�j`"�9�-`JR2n-�{�^�3L����`�\c��)�<$ ���3���n��.���5
��甙�r���%�S�4�cm:a�ԈT�iX�Ȍ/�}�f�������Ĭd$.kA ��$����o���#�n��ō0_�����3j�E{v,F�o�#���ёT��_h�>>L�6���ϊ��|v�}��<�,���{���(?�M�s}<Wv���l`��0!��v��;S\XJW�7�O�&A�>����RT+<A�
�ks0��1~1ɿO&��NV�@kU����^�a�Vl*���I@@` ���Q }y����L__��jxʾ�!��ɔ�WLտr�P�F�1�f��_1��mmlm~H>�E7�@�����$N���U�R�z����_Ljx]�����n���,�]��ʌ�J����쏙�u�Aj�*}x:"ڪu�!/��f�E@ xdh����:2��d� N��!k)����(��������}ˀ�;�w�����M���iy�c]��u_��	�ps��f���w�X���[����%�v��S��ұuT����2$�@�#0]ȹ)㣄|�&b������_���=�~G��0��+!q����{o��q�sӏ$��^�R�?J������,e�Q�T&�6+���l8��`��8l7�:W�l�ً������QM��s�@�uٺ�@}�x~umF�g}�j]P؇	n8ccbV;�v��՝�y�n_��]�Jd+�_�������KC�<,n�[߷9D��X!�B�����NK�*׀Er�y�a���ק j!q�RW�m��-O� ���ei�[�QeM"��?�U\{�����8{g������F3��@	<~<+�����?��"���ׯ�q���4d>��dRZoMܖ���t�������+_�ȿ��J���i�'v��|��<��	�E��6#`�W������D��P�e?�#�Q�f{
���w6K׏�/S/=�~��~3_�*0bM�&2k���ޞ߃�V/��"����`J�ӡX�(cN2_5&C�.�`�<<N@n*���L�=�
Č�1p�h�E�h^ݼ7Z0t*	?os�Ng��G��<��4�����I�cX�����T���3Ѽ����5@�W�"�l�Գ���ɢfϖ�xq9�ӖŰ��N�l-kO'_ ż�k�[��"U�m4��N�X��u�a������| ��(��׾�8յX�aB�G?0�$/�>�涷�&+���C���dD�T���L��c�{���@H�;]R�@��^qj�=4U:�h5�_�������g�4됅v.J������� ��o��o��#a���.��(�����b���#wgj��O�wV�⤜S��e2K[�]�`�7��a�1sZe��1g�۹&���{�)f�N|�jy����"��G^}���b3����&���C�^��lDa8k��**W�|��ު�@�`�&҉83T�k�e�,B��k=ֆFF������6F�����Ͽ��T�Ԁ���A=Y��6���o��@
��C���Gñ+·pN��8ʔ��<�_0i{w��*��㞾�!u��/�>{)���1�T��u��rrU��DU�t��wr~Θ�f����x&�{g��C�O�b�
2@?�J�0N�A�X�^��s��O�]����S��.g����*��������h��B�Y�vv�O_T��;�i������B����0R�I[�o�#C3���0�ɚ�l��n^��5�G8����8콜N���?�P��,�}�������ڸq��L�3ȻW�d�x�)�h犄���#�IDC͠�k���r��jkO� �fEt��6HU��x�M�����exl��3Д��R�@�[�a��l�-Fƌ�q��6�kHZ�s�$����l2+jXntW��n�g�da�c���	]���X��5Ԝ�NE9��s�v���6�o�(�f�x� )�O2--q��ޞӲSS����ɗd9w��7#���UK:���*��7���$����/7a�:d�Q#=u���\o�𴇦<(�щ��,OO��<�=%ȯP�;����:.ʠk�niIi�AB������{�ni	A@��K$V��������y���ta���9W̜33͹�W#֞9N[&����*E��@�8�X��Z��7%j�(+������a��ʸd`n	�̓(����nB��`|>��N��u+q{�3UR4�Õ��%�9�J�x����%!�^<�:lK�?x���(����!�� f�r��:,����o�mn��f�g���D��_�A#bQD��N7���i�y��������x�:�����b%i dzr2Pq�^c�Zf�?����Y���7|�ݩ�/����
�mk�S�þ��}!Q�*of�e�?�P@��~C�E�tۡu��E6�;	�k!j���8�ߧ���Q�g[|��!(�ZA�������s�,�w6��& ������Q����iBޗ?���~<˼��Aq� EV}0�
.�[��<���y$y��Ǿ:�#0(���� ����x�L �l~,4���?�B�bp�N���8@1���-u���5C��/0z^$O�T^�nL�o����n���E(E�����!��	���S/����}l��H���ն�☒�Η�R�N�a�WK�܁���?7�}������#����d&S�)?�,^;�0��#iC��}Y��uI/�efrF���N�NK�R7Y�l����Y^w��@����CQDm� K�6=(>[[�V��y�nӒ�h+�_�8��Ugh$�;��r � ����]9���n�����'[�_��|��U�9z1�V.�$r8p1@z��{���f�E�R��+����;�����\��lV���FxQvpH���P�V(�X��B*cGk!JW:NOU�
-�����n��?���l��Zv�R�E��%:N� �G�>�[�N������O222��b�q����
�X��ܪ�R�?��Y�
�O�ex�Q���^�3Í��\��텼��oSi�ؘ3+��)#f|�\���ڇ��,3����ղ�QbT#��@������N����AV\ύ�����Qdvf`�7�33�`7w�f�~��`���"ٳ#zE�o#�Edp��n����i师.՛�,��yu���0w��/1EhH�'�MU{B�(�<#>=w��N=����^}w	Xj��)�m�!�f�7g��~�u3�U���gY"}���U !�Tmo�>�^�{�G"ܔ鹲�p���	Q�7��I8�R�G��\��NͿ����\������"��ÿjh�ѕ��rH���vԶN!,v��������A��
��9)���.$��@h3G?AO�����2̗9[)S��c;�{!���B0,D��$���w��-�<p���`��`?�`�Mr� ҴA(G�[G�f��i��Q�vE�N��&ť�ϝSߟ{�JU6�I<� ,�Q{ɢ�,��!"̍lZX�T���ݵ�j$nVD��dLT��10e�뢐ب�pī0��_��ȳ�4���fs��&�قT��dҊ��w �G���8Hf��:�A��7sK{�F �	Ʒ�WF��M\K�Qw)A�[qB&:���v�_ld�/��Ǝ'�x�� ���u����C^ڶ(-�� rW7�r;��S��G;�#�B����DDD]��J5WaL1�cT6Z���(=M祒�e���O�cwW��P��?���q����?/�����-�����V/�fcSȊl�逩����S>�����S0�V�� +���`�q#h��o���/06��خ~�l��4H":�@x�T��K�Ѐ����ג�f� ����f�0M�}	�,nٟ�PЏ��(�����X��o�p7ѧ�P����l8�a�x1�J,���v��	�=X��Ђv��L��)����p�KFFb|�F�$���a�j�;��I�9�!qC�\۸�Qs�	[]���3�u��s�Wy��3�|���2�����s�TO�U5)���,��E��<K� �Aؕ?�&���Bq���.
pP��� ���܌>>��B�M�AE�=]�����5�
�vFʘ'ˌ��oO���¢�<�WH�VOFU��D
�
��j��\�u�Ӻ����yk1vRABj�����m��:i��2�`��j���dz_�ت��ֹ����3���ߦ|��:�r��Zcqq�)�n���?!V��M���{J(}ӭ4e�5��m�Jղ+&�,�0`H���/者<7��Z�}�0)Qۋ=���+Uc�����n>�#�6�_�tD<ś3S��#z��2�p�c��·���ד ��I9g���+���a�J�Ah���D3�7_RJ�lgJރ�S7mo�EUII�_q��
���Օ3#c@�Z��]�/b+/<�4i�X̢XSo��h�k�'�*7�Dȣ2�oZ~g���:���&��1�x��j���b���h��%�g� �5��K~[�K�G?��_KI�۬��UQ�^M�fO����f6S�&�]$��C3a�Y��{榛�}2�Eo�M0��=�a�[R:� ��dT/������l���;_?�"-�jN2��������E*l�CJF&�m-���K�Q�0ѫ�3�æ��#�TUUS��e�,~�9������x��#N���봨D/켅�|웜������&6܈��
�ML�G���>�і����T�>�Fq�z؛*ӂ�΅�K�#c}���TaOT���m��K57��$���̛���t���&��y���܁9䚨��ihW�̢���b��~����!s���I�Pr�uj���<�U��g�V�#�D��w�T��=�Vu�GC =P��pbLY3��h��,S���#lT{J,�X��%�����Ma҄�-ɖ�Ӧ+�+3��|�$՟����M�B�Exi��}4*#���d`�ZUr񦣤bs����馘�� ����K^n�����-ڈ�A �S�.���I2�3(�����loۯ��g}�.���NP׿�Y�"�����84�w�o0�"/�j���$���&���-$ue��67=���0���Wg6���e��|p�5�a�p_>f&�Wh�R,UM�X�f�cM'Erp��F��am�Г��A�XiqsíF���Ja<T��p|�T��fC]�~wU?aͮO��l����z�*���%j��hF�>~����ى,q���+��Ϗ��a�gXCf3�!�/��e~9�Dr��ˊ�D���J���M.�p�V�������α��(���3�1I�3�h�1�K]CC��3�ml��뛚���������*1C�T��s�q=�r��Ih�c� ivf����~�B����gl^�]pj*���Č��ۼ?Z�T�W��1�׽|��5��W]_Wq��������Ō����X �:<��˛*a�ozL��L�_2��fL�+ھ�Vv3f �yByjj�2+�錴:FΚ��t���|�}TXs���kǤۨ��<pf�[[0i#�/�P�8����|��o�\����Km919򨃮����-]���� 0�i<	��!yV���E-�/�H �����`�M��
�1��r��C�:q�mV����2�4QO�tś�v�\o��L���]肂.
�Iw��*�	K��S�ݒ�\jR������4��c�mK��K��>����$tY\z�jl��uX/�-HW��u���z(eнѾ�${�� z4+���II�@O�yt�GCdf�f�����º'�V��.$��w1]p��k��h/!���.C7�m��J�FO��^���G2�	�	�#�x����"�M����%+#�'���r���e�=7Vu�2B�4+�y���|�F-�X�E�"��B��d6E-�y�����u��F[�8 h{��7�~�J���E�P��sr�(��"�X6����bw��= ��F.�`���	/��[9���J����[tt�-������}w��B���li����,�ͥ�E��=��5�>Y�nM�X6��C��\B�D�udL�&�D�)F2_�-+d�����-��	<`Nm�ǲ���%8��2�;vgׯ./�g��xy��-)�d��q�{E�A��}-|b5y[�����CG��pi�rh�T�$96$N�@1�ⷚt8G�w㣢e3mWo2�+�/I0ȣʲ��̳=qmmm�k��+��S����z�	!��i\Ɨ��O�4�)"��&����-&
=�8�����(�5�)�o�X�b.T:��i��(C@��ՙ���u�E�Em�4�m���a��T�:<�܊��4�b���b�JJ:q&�E�F"	b�v�+U���J7o�:�|Ӓf��뭡�̈́���B�mY�[.�ށR[��'�Ч+ ��ɠ�Aɵ�~�\ta��H'7#��l*�Ŗ��
�� ���ύ�O~��Jc��vT.]&����M������o�FO�D�e��ߛ6��=�u�[~��=(	���-ӡ^�vm*Y��\ڟ\�i5�����'S��܆aooo,~�C>@ �}�øV�I:]y�f�1'�RrہֳO�p/d5+T���s��r����c��L��k��|o�I2��A���4wr����f��7?�ё���	�O������̜�֓?��;�M\g��a���ō�WhGL�(��I�Z�9�x��[~�vE2����O	U�B�� '��ٶ�ːP�֘�Y�?7y��r�(�ڻǬZQ"/\���?�h�Uk%�ufdf���A���A�ma��j���Aј�8]��z����~wz�O�M�!�w��o�	���"**(�&��:&��%7wp���l�����440"u�������0C��*.��B���ƥ��D�<lh�I��;U���ҋ�Zo/o��A@�Z	��G/�Y�ɞ����-���]��-7�U4g��b����/�5c��:�D�Q?)۸���oB��c�K�����$����	æ����D} &�x���6��3��v��_lҁu9H���B})����]1��©au��}:C��&�&�e��$ųM�'&'��L�ց��V�b��oqA�f;���0S�t,s������韛���VC�����:@����7�|��|�u�/Q`$�X��R.t��b�w�D�T�V��+E�*[�G/̚ϣ 9����sٙ������6E��`yl�u��S��}��D�_dE2??<���<:0Ak�#�����1_:GA:^��d�������N}s�ˋ'�ty5����0cb��`��Ľ�:N2Z</�zrv��E��㱔�	����Q�v�y��ďV��Ź�c�R�pq�\t��v�eMK"Xa�|�� lެ7��d%��wT#�CrֲG1b�8�`�����-�ջ�1�5Ir3�������f�SՅ�$�7y�	dC��f�Z/���m=n)�L���;���r�>v�����f*�g>��C�R�W*7��H`+��n��b�
��b�E����\w�����i]8���+L�i(4�T,<6�T��8,vrwg��y�)��qP��y��GG�]\�ĩ��o�./��D΅O �������St�y_����7���-$1[��H�-@]e�c�ߏ�^L2?���!7:\�S�h�Cj�mx�3Ĩf���q-��R;�f͙*�:UB�}[��gm��e�4t+�WX^��	��>0˩c��fJ-F��my�l�!M�脬22u<�z��3y0���?111�U݂%����E����/b�s�6�(h�ȼ�҇�r��p-z�+?DJR���`�0��P���Pc-��zjVf;ǹ�}�ޤ����W���i��ߨ��up0�(�[�K���dJ�Ƒ�*���)�]��D��툹���͘f3hD��̆���P�p�Z�x^���Y'!
B���n-Q���4B@��^�NՅה��"_~�������F=�������8�M���Z
񯕕�	�zz}�~��<�l��q1KR�J���z�;�Z b�C��:Uc]c���)B�:�Q[�i@<�����Qsf��꘻��;w�vn4|�M��Lu�<��3�^v�go��B2C<L���`�;���c��Pj'�8�����%��S�-������D�t��6�������֏W@B���s)()}������Z��5�C��7�^d-����'�L��Qe�9E��d�P����N��ݽ��d8a��q=�강͏�:p�ϩ=n��B�x�������-I�4����x)f}0�@�U��oTC��y�r0;���x&2��.�Y����f|��g��S�χ�#�m�ޠ֗�r����iKE>ߓw�������آH��s����c�ڪ������N�a����e6����9�����G�Un-��(1"�p��snS�x;w�2�U8�6�}��޻�f����vo�f�y�Z0ڥ�Ѷe*j���f��Խ3�B_�����{<=\Ac�J�p�"v�Ј`C�Hu��$�+>���fs6�N��.��m>sپO�w�[JI�'������!1qW:�MKh����BU��ƣ���O�^,�'s��_?V"���X��6K��M��G��l�I�!1 >M�����p�pꏹ9�ǋ��9�%"Y���c�_���d�}[۷j�VaL�t��L�.cm�Z�Z��Q������]h����_%��^�����ۤ�QUU�S�� $������q�ۻ;��A@��}%�A1�iA�<rX�oqJ)�]�V*Y�L�ܷ�_ǁ�W��+v�_)1!���F�K*�?5-��"�[,*�K���FG��Q�ՠ��2����E�ϒ������܅W&����ִ���m\������ￆ��5��Z�"���Ͱt^j�_h������a����6��ʣ�O��JK��,G��Xg,08z�G���:RU?d�	n=�L�Z���!S|��ZC��!�ښ�w��
����D��֨��κ�Yڋ��ۓص�Eiq�G��X��pv��I*}ܽM�Z�rh�WFU�f(N�\r��:�c���8ߜ�>�X�g^� ��_����h)r��f��i �i�yt}��l2�ܪ�̹�B����դTѱ�u� ��J	.��� cLA�H7�M��B��嵉�IQ=a�nr��,�H$^D6�.�	��Pf��h�y������z=�:w��S;�w�~,N䱉�^_AQ1}D޷8D�þ�60,S�4��~���R^!E%� _���C�7��o�ܤ�b�Wq�����U^� Y �,�ￖ�9]��
�A�˧�@O ��D�&r��9����p��;���n������X\��8����@��燐N��=��@�zďZ�J�[�A|n�HN\���@��8���I,>O���vJ&Z�X�I��=��7/�(9��'o�gN�׍%�Q�G�_]���uT�~|�'���Ϗ\^^��bv6�勛��w����HiY��J���*��PAK aA	�cJ�����(�� �$���2$�/�`H�緵���L�X~=�	���; ����ē�c�8.+_���9�G�&[ȣ�S�h���m��׋�x)�����.��UN<o`p�LZ96	oD���̜�;��{u����v�.UI�!v9�A�����D�,7x\�Y��2� ���f3[�ǪD�{x����_�����>#����/A\�����.���O �"E/��ˍ���*�W_{�GT���f(�������:cJ<��֪e+$�,�ZD��.�Ӊ�Nz�qq����0����%;c<�O-@�~e�c���=���A�]Ψ9��M�n���{e��p�&7�����>��U����~�j����%z��].=;۬�L�*AԾ�s2S�����~��9�awʉ?G��"??'��ѷ��X�]�-���_A��o3��W�.e)		��W|kC&���m���f��xr>]|Xă��=��2ŬO���+ǰ�L�RT-�e����	��lN�e<q�SSS{���e����
s�����7�L�jtt���.�;d�7U�U���}}$	�G�+��2�K�['r3b9�o�Æ�v=?�AG��]�+_Z�wAإJ@!�>�@�|�y���?S�9���L�s/%]ќH�B�-���"��0�\�t�h�%�'xb�_�j\����~Kl���:Jء�n����b���ڻ�?����~ ���;�d@�O�5�D��Ӊ��b��H��N����?:��Q��(J���0��LU���S� 
��=ٹSd��qJճZe2
xQ O�A]���v�M�)\C��G8$<��Ǻ~V..���Ο�C�LU�nTs3��b��F	�b/�yq0��Zfg���y�m)�EQ�Pޓ�I#��H ��V����\�ƈ�����v\ ���np�����ˮ7O܄���kik�QMOO�R���]�ʲ���w9 M�a����w��������3Rѧ����a�<��@��G���R>v�$1�+���g�^�]�D���S��}��
��(�\��Q�������&i���O8 §N.ܝ�V�zl�]E�Lx?S!-:y�.��P�9���(�G3�=.1ymaȂ2QQ�̄��>���!���rڪ]��W���BΒ?HѶB/*�h�!i��"�Яy��FSW������24���%u�#IC�\������I/vp��T�p��-���}A���soh�'�ӗ���_��59������z#�[�P���1�y�)��^a�=ӯ�v�G�ѐ�:���yP���i�b��{��ə7 ޘ(U ����;��ݢ��$���m���p���OSN��Dm!M8ddc���]�#i��c�[��aW����f*���r܋\{�O���SUK#��&G��9G�	080/�R��0�vpAEy�B�3l������Pu��/���WS�+�ej��]�`Q\�X*֊�	0B侇�s��L��s-����,������ /M~w�>�^��i��ݕ��t9 M�de�]T[XXp P}S��	٠��r���G��O	cd;��&7�г� �7и�(�u�_ʌ�v��ĳ�fnm��n�H��.�<宒��L~��;��������A�'\�W冭n/�7�$ဨ�񃀑 3Y�=�*Afe�>T�+�����bx<�s��ȶ����HICt�r��� �\|�kb3|ťh��m\�����WXI��
�.A�A�K��1��j:�Ԩ^Y<!R�*�C[�S�4ih�6��@��|�܀L��}bUz���!c�W���I[\�V��M�K�j�|�h�oA�>�L�����)靁 �Sc ���#�>����2y�3�;/�;�v&�]��)^ZڅMW���I��<~{2�i��,ysU�1�+� =��v���QG`�ķTu�G6��uf�b�@�M>��Y�2�疵�3��A���J�Gq$��YS�]�j�]��J5h ^��d���\Cp��)Ň�E���.�@	��%|r�l1&�N��Ï�B-�?J�.�m4-ol$â�3R�q��{Ϥv:m�����b�,�mX����\�PA I��K�d��`�%޸�U��6�`������F�쫵��n#Z�#���|tZ�BS�S�T��Z�l�}F���׮�dac�s+��o~��z�5�j�L�A������?�,��rkl0ᾙ�OʢQt�p4���۫&"_pƘ>�atlYE��Fg���Fլ����,|���\h�S���fI��k\W�����/�7��P�N�)��`p�����0ɂ�lB�U\m��������ؘ�+�p�>_��9�)��	�K��)A��(��d��_ul0ZR�K�X����7'I1��Dk�S�zK�?.�V��9;t
}3�<Dk��*��t�J($��X��%'*���m$
�N����.@|w�b^ �omi�����s1T&����y���3�!��I^n�0k\�uX���`:??7m�䒣s�����G�J���E�0T�5�J��nRM�w��8�����������ձ\��i��U���Ao/����JIF5�-B����.��q�zÂ����%ݺ����ِ�t a�ĩL�o��o���� _�½!��2)��������᎒�(�vL)���Gi���r�[�������������������������	���6Ϸ:::�K�l�Th��Ri�Ir����bœ��1�����Qs]�Y�8%���<�߰���qPJ�(%9u^��y��\y��S1�)�'Ա�8��q�}�r��$�L ?= ���T#ן�J�<D9l)	H�i�oArf��t�\�K���
��X'����~gN����f�vT�������͝WZ*��*)O#�3ʻ�7�G��ZDD��Ieǅ�`���6~�<`K������L��N2�hs�I�?������	}�&���1F�u�t�(��B�x��0���J��r��0�,���K�K�.�������|�ikm����ؐ݌/�
��%�6�]��kE�4�Mn5"�Q��;x�(�pVT����"����p��j.�ـ�I\����E��L��F�k��o0WO^>��F�H^��#y��cj�c;:==���Y����\���l�w~�%'?���E�FEú4D�I�w��Z�/.�,9�$�+M��ҁ S<A-�Oq-�1���(
Ó��T�@�	����#/���Dc0��S�����uGlׅx�B�xm`�'��O�-zP����H���^O�A��g�j�,�Ᾱ�y�q��_t6�u?�������/ZX/)�|��]·܌��㝚o0�*x�85[MB��	C��5t}�}�^��E���C��R�����gx��۔�S$�vke��U�pÜiH�/�p��滴	gW\շ�d�t�Jqr�|����C�8�ˢ�{�+��9�Avm��ܼ����R蓉�h��]t���w�G��V������ �#YF�C�}��շ�9?t��m�p�u����)���ȱ�}��?�ތ��Ye1N�����t��r����Ȉ��ac1$�nD�C������n�dp��}@o�ˀ�3bi�l�f�:�O�'�[�Q#l�Y)��3��Z����fU�=��c�v9�M9�c��3G�)��n�� ���GIR]���C���Ӄq&��5,ދi����nh�0f��ix�F�M�lɕ__���>�rI죲�z�Df�%W��Y�퍩�@ <rMK~@>9yh>3&g��̓_�v������G� ��K�,<|;䀒]�{|�k&B ~�
Md0[��_�_O+h0�L̹�� ߅c�+���p���c��Z�}Me�⃛@�O0�3�~��4�C,�׿�䦶���c����]�~!@�3NK�X���J��)�_	y�!)��Ī1��W~���/Ȟ� ����V���j/0w�������*g�]�:��!�'�g�f
D�O��@)~������ҙ\Z�U�Y����Y8&���U7���@+*x�ٵ��
Zp��v=n�������z��\���Qe�^��j�FFF��M�� ���Us6M���ʚ�i�Ӹc|���63��s?t�|}|W�.#�sێ?���)k�..8G���X�G�c�[�{��v|���������F)"B���ji9��*�R�^�i�D��f3��KȮ��MMMʹ�%d`p�`D~@�|(s��+s�tY�!U�SK�,	�JB.M�^�1/\ɲI(V����d��:Æ��ga�pʭ���xm>@"UU9x�
��lTҧ���@ Z����066��v!{sjEW���������/������5սXRr�F)+; ���m���o+�t3��J�b ������H��0|��ȓ�R`b�0j.?{��^RQ1��L9��/�u���!��駵	ؤ�pl{&�[A�ӟd��JM��z����{��f�-�/��6&���5�=l\��>�ᑭ�k׌CLl��ğ�_:�k`@�vA- �������N(XvD6-��?�&v�+����G{Ͻ������,�w��KN���nnnK+�@���zWW�l��v�8��Xh�uh]�*�2�"qܙ�LNI1�727G�k�&u�2���jY��!���)hS���߮,�%��p%��J�:�;��������R�κ�hV�v�1�1�ې{��`��7-�Q�R�a.)���)-m���w��ܔ-��]��>[JTmd"���[&��ʊ��̻��.�bE�k�#��0�#���8�����U�X`9�7U�E������f�I:��~�Yޒ�lb�iT���T�%W��]t=q%��ף]��$e��E�rL��ih����d���}*I��[]]�,b����j__S���7��}��'y�Ғ�䗕Y����O	�G�jz/0h�Kݢ�w�n&�l;M��~���[�8�[�f��ʋ�#�ذ�?�xy%w4�t>��A�*���� a����'|ԲϚ�l�;�-�_�F�s��f�R�P-��-%�7d	�̈́�Bƙ�(i!�;I��="��m��8и6��(�h@s�`EV�"+���)��mg���p%�k��r*}���
�J���;<䆛�i�M� ��~��O"ek�{�4����qQ���
s0�(ÞF0�A---�1�\i��{MY?EC�b��ݾ�?����3痗t�ud�S+��}j���\h0��>�����_6�C�໿�1<u&$$, #�P�����ֶ_�wQ�{t���X~I��qi���, �#��;�I1��}��y*!4n�0Ѯ\����ͯ��&*���PC�goo���頦��S7ڴ,i))�O\��@���Ҳ`�.�$F����띹�����{��dzlC�_��s�&.����Mq�jCb���	�\[�"�9�R���ӵ��&���2W/ߡ5'mr(( ;��K,��y{��g�cm��6;����)L3��~���k{^��E;��J2T�#��Կ`H�$"�^��vGp��ow
V�F��1�j���_���nT)o��3 �'w��C?��].��	p:���+z�������3�#��������"�	�i��v� ݠ���s-�:�sq_�L3T:{C���_m��3TӶ��40����6�� \@d$��{~Gy&���C��{Se��4O%����#�?�`��}��f*f�!:I�Z�}���鸊�摑��<ZT��G@ �6;��2?��i�M��kl\%�X>6d�l���t�8"+ЩjX��/ �V�)�\��q�o�o&{Δ��h��N����_v��<?���׿�i�<�M6�;���;�\NX��_��PٳZ�[��hJ�M�e�¦
7�;�2vh흰#�L�K8tJJ�]M0�{���Od���u���e����dƄquqYI�ȑݿa&@ H�OL[~>�B���o��B�!��8��e����h�J���)�N��K�灶���StT4���:��aj��9!��*�6�{	Aw�32H`D_c���9��:���j\�l:5W����(�N��n��qGGG�����+�B�b{' g��3��a��#�^�B�����@��o>�ЃζF�*�x2�xE����=�#�����x} ơY��,���uV|��	嵔
���6�NA��N�?�gy�������i� ξ0���eA�v�����W�O��/xQV��A���>"�=p:��
	��y�)?�(ι鮭��C����!����3�~�X����֯���רڽD&R3�hMI��>�»�y��v�o�9�V'�ҔeD�|���4�&K���3�l>�nGwG?��ĸHa�� �O�� ��־7B�s"�1�,R�"�G�77��F�B>���4�����fx��� I���&w����`�_k�gj�۽�tFPPw���`��Ǐ��_���|}}��)�����o���>�V��3�Q����.�?U���q�R99�Ţ�M�6�%P�n�+����,--�N��![�N�?�ᶺ�t>��񅆅�` ��ͨ��{��i�{PaЦgsɡȎ����z#�&+e�L�ˤ��F����۱���ܥ���_���8��J͈��+�6�����O�����un���G;���<���0�)��U'ſ�"���n,�xA�h���P$�i����b�SC�]d���V��qP$��9l�;Ƞ�Iæ?��O��p����rr%�������^a�t��BGZ�N��^��L��f:.��e���0��L%lC�J@1�Vj��Nuai�Z^n��܎w�!���Κ�?0Z�u�@�.���.���g!R�3Qǝ�Ke:,��5^:��$��(�Q��F؆O�3����l]G��oyV�[ZH�� nN�`-��\lu/���'�f�I���Z����������N�7}���B��R)��s�t��#��v]b����N,?�����c�:�g0�%0��Gb�u�п�ͭ~��ը�L�S9C|���pv��Q}\�\Pw��]`A�wS48�giJ:M�b'�N_#�׷ۂ�1��L��U���� ���g�u�Lf���Ps�#C���n�BLlƙ��[��P��g�zs&��z�Y�[#�H���B*ŨF��Q�|�c;We�r���DO�Cy��x3H#+������AЎTT\L)�t�5Hԛʢ�0��8��<)�`���Z=:Y\RR0���jR�� ��ړ�U����Z�sK��`�x�!Z��ëI�Sv�uz��rp���J0�X�W���WVQ���� �-̆SPZ�V^^�Ns�1�l` ��O�*A
�M��b�}�ƈ�^�����ӏ�Ŀ&J�䇼
/�E�L%@Ps��4~VBP�pu�����3���Rl��u���]���r��0E?�m�JǑc%4mo�r�}3��^��e�A�[�E�+��W�#̼����J�d~�k��/��������H�X� P=r s0�yUU�ִ)������ɨ	��9wT����]GHII)�&�y=AE�!�ٚ/'�"d�P�[��n���vZ�0�0]�)^e��}�hAA�5tY^����1�wU�����ZX�pq�����|�k;�*ho�����fNV|4�T	��B'��ZS<`�u�Q�x�t�&�+�4ц�x\#��/����^��zкR�d^s3ߪ�����3G���,�Zr"$(d����xe����5���^�݊S3n���Am+&�[sM�19"�}�� �!���e�/�C���Zx�/����М��ta܇1��{������ �CCyH����;lH8-2q��u��
���[m)]b�)���Q����M ���#P2�#Q�wك68��D�ϥ���*	���_C�д���[j �y_WW�5/�x�@dR��b��� �}_y�R�OG8=tt,LL����כ����I���p$���i�a#���P^!���Ғ� ��_�2��`^�А&�-f�ｽ.��+筕�T��-MbM�L���KY[3�2w�H�A�ϕf'ҫ;�� ��M��l�wo ����o}�Z�X�G�tv
z���H��ʀ�O4�h��T�� ҌG%�r*c�ܼ��RRRo��GG�Vj\�z�ׇ`n�6�n�`�k����, h[T�xlqNk��g�����{�4���!wB��y�!�0R~�Fy�}@`(q��G���3A�lNK�����Lhh��g}�đ_�S�11��?WR5�i=??�,WD�:�uO9��;��D��a��:�̹H�O��!��H�b`��H��(�@lu�Ȳ꛷�kk�K���ͻy:�ㆇe�45-�[�9���޼��g��q��r�.����������$����w�W�<�_�*��
ev�0����b�'��� e<�[��w�ᠷu���`@����@����\baV�lmYܠ�R3�%��#ha��ֺ/�������	^�G!��	Y�l����D�;~�_�i��\�#���� ��qeM�q�Ր-�K��ph�>�T���v��p"D�����e���}1�*zm59�@X [��AS(Xm���J���*�.��tl��]�5�n;͗x��y	Ŀ<`l��#�e) G;�2!=8�D�0�8ർ����q�ߎ�p^�R:�T�����d�x���h�kE:pa���L��q��� ~z���D��'*�?��ħ'CJ;s�O����َ�ڈ�J�m5�I\~�k����Y�&�<�q����VT�,
�h���[�Ǝ�!��ss��\o[��u.����2�һ�P2��ޜ%�7!�+ �����GW�KjqM��6A��^o�|)Y`m�i
�a�L����V�M�0 i������X��{�0�K M�LsqEN��l?�9y�����n&wn[�@��
�wKa �������V��O#��\���4�leV;������<�D�����y�F�[6QYS3���q�>
V>l�C�N�����Q��Dr��i��7yqԂoë�;�����z,,,��a����l�g�^%� ����GG��z7�J�����r�/H5��QM0�Zɀ駪�:�!�;�708�D��4^�,�K�J�i>���J����+ʹ�3��3��KM.�������hZ�0��/Y���zvzG���Hچ����ԟHql'>���ڒ���^^^�a�ܳJ�����ӗR*������zuQ'�W|�3�wU&:_�%^����|�vT��.�;m ��a��_��er)g�nnnZ�ۇ-�rv����e��l"���m��^ER��(�$�(���jG���hY�Tn8��B7�w��]z����Λ��t,@����Ay��·i3k�ɟg�Э�f�~ �e�d��,Qy���.�e���n�Ly0@��]��:�Ȫ�:%.Z`��t��&щ3M/(�b���1��;)����E�d�D��e��F�V��{`~�̈��G��f��s���_�*#�q�n�m/����lbܦ�iAT��y~yG\��]R���\���5� �;�ٿ�o��� :�fhiҰWf��K�vvf�ZP�kb8��vH>�]��0��4l��-=�HNM��T�<K��p�3��i7�S��1~�w�[��`�cx�0��"��>C���-��U����QM|���4�WB��~I"gM�;��n\�S�~����
�8�����m��\��C� !H������-x���{��5����������֚E��g���ޟTUW�����-;44PSS3q0�t��:jv�Ò����r�1؆���I�oi3��Ʋ !�Z�2"8��>hll,hg�����p���G�����Z�AQ����Ϸ�T<8��}�P�1=��&(x��r�{�u�MC�>Q���)����XYm}�e��״��`� ����l=�H��m�7{��_bp��C�A��x� �tS�׍b?r��5V���-�Z_(�Z#�}�5��9�$M��h>�+�L�)yN]���l~$�YmT��T��+հ1?@p��
o�g��M�
O���|������s������QdT���~����ݐ�g�=BL�.�~}�C�Ռͫ��0Ǡ̌�͕����rK3�66J� �
��cM\�Q�,G�oH>Ȑ#���#e�D��̬ۨ���@�Ȅ�q=�5P�!�)�p���8�;�6�k�!�oM���r��$54p���S|�ڛ�����f�SH1�:D{ �[�t��Y��u���Q�e����c�����vij+�Cc�wT>�bi�VZ*5}��;�C�RI�!S���_,��𚆧��4�@��UȠ�����*�l E:ͯ�aŃ�u��ʴ`�蠸���m���ƒj�����qg͉���0"�g%�S��?E�ި�2i!��Tٮ
/9��~��S��ښ��8�Dc�_4�w�E�4�A��+ǃ�g�ப�an�;�L�$��d��r����+H/֢m�.'�$��	dn��ݽ������v�����XT �P�A�r��}�֯ϴ
bk��*���*GT� E��ߐ�~5�i?O��������r�0c�tȞ/@<�RR���0O�9}�����|��#J�ғ�+�TP+�z���)M>���T�}���#i����_s$��Z�i �d�uT7�-E &�m?�"�V����(�?<�~�|��mp�%<�^��^x'� c�C�|KY����>&
B��Lq�Kʤ����#�/�����Y�9�4Quuu�22T�G
�߾��5Z\L��@;�m���-��I�+""�$*��B z��Lq`���냺�7����&�2O?�p����L����o%I�:I��Â�"�Gl{�+3��i��CzPQQ�u�E����*Z����&���Ĝ�8����\/G�'�0{�����y͔�D��a�	���T��}������_����a��<����H37 Juk��.gזe�ۻس�+ͪ4!4v�PǸ3������.T5ӟ\会,	���v�V	�rܯlǦ�������h�G�ϳE*5_.���Z����� ��u��hB��3���?� ��k5����*��?d����L�Ĉ��Wu�S̻�>(�/=T�pM���T ��\^��j��{��Nvmj~K��~���~b[]��ݰ�#�����fN\���I�6a%���UQ��k�ֲ �j�o~�{߄����1�ɫ$J	�%vy�J���i2�tu�QT�������o�]7�uv���s�r���gl�������]�����xb�珨���:�ٝO3<~z$^a�Rmil�n�1�Ǚ�u�c�e"-m�G���	�⧻�l��U�5s}�fk�9�� ��~�8�����Si��F577�D�Y�	�߽�0�덭*��t��_�*����S��C5���bRܥ0!���Fi<:���9�����+�1��2��͢dj|��)ͤf���l�f Gd��r�>����L�F��'o~g�=[�c�I���!�zx���п��^[_'����XxHϵ����2���ľo���ZҺ����m߿O��Rݾ�c̺\U�вg�����|jHf� ���ed*�ǺjQ]���'�q*��`��RQ�#d����p���#��# ��ZZ����muF9��P4���YX�MLh�N��u�YYY��_o4�لS&E�^)p0�l����N�ò��8��S�kd��d��}{���쵁���*�u���F���Ʃ�;2�#`B?7w
N���QS	))8@#:R���|i�Q��o�|�)�O�~u�_Ad�x'��`�r�Ntr"lY��L�(7@�b�"Rh})�C���FDn,����ov��w�|p�ܲ�.:��?�"9��a!5��=�������<����U�o���m�M&�zeee*0���,�,��]ʊ�xQ�#���Br�x�_罦f�,uB������R���G���='CCCʽ��l���H;��!�4 ?W{佉;T����>�l�m����Bmm�ݖ
��Q�Jݽn����ۊ{ɮ�o=�� �O�Q��u��6$�v���o���xI~,EҺ�Cv�\^�njj
Z��<�Wڽy�����5?�U�� ��yF�膑V�;��\�Y����7^����~qt����kY�Oՙ���+H���"Z�`H�2�MHL� ��楖X��*��5a���Y�0L@�c��.�YP�x����\�D�֯��|F��|�(�U9�o�f]R�pg-�M�~ �1��!PYl�������}°kj���� ��ų+I�`L�8��C�5��f���c��t����g@(��ңM/���uI�������R��H ����M2Nv��}�ڌƧ��ϣ���ʫ�@����"}������2���ީ
i�´�a|�=�Z� 9���oafX9d��LI,����f;�K�����ǛM���*{q�9 =���xnoh�s����QS���D¢�"zF��R���H�U�iEm\���O��G?f됿;���$�xY��b~O:i�AG���|ú��{���4�x�Ȼ��q��U�0.A��Nm���}}}��=sɟsé� ena� HU�������}�i�يͱ�l��>�9-н��3�B��w��+	�eb(�{XuA\�v�92��3�0�~Jɢof�t���Y�v<����	�Z��sm1�qT����eͥ��l�(.���ێ�����n��*���T;�b�''gѹ��+�f�gƷ��.��}�frb�GYU5�ʌwO�]����z1*<..�+����o޼�������l%Ad ��Ʃ�U��c�F?��@��}�=���W��|�5=a#�����91�����V�J^r[W�����Mdi=A����'" +����f``���� ��j���x.�V���*���>G���A���{l�X��nǔ�qV�c�t�3|i�S�w<�S��-C�ܲm$G�������5׮�!9�6=�$��:��.}Quu���2LTxv!�h 3�&�L��p21IjiB�i�0K�ަ����/�jO8���R�{�� }����-�e�BS����°�$q3v�BEJ����C݌)α�;Y@:�tGRM�`��p����y�s�5(&�%(urZ�qd�/5�" ���h+�Ã8ν�=��B}�L��8��<	�m���B�wz��f��pr�в��@��[��͛���n 9]\��b���C7d?�83/���E���׸�[.�l���������5)�otD�a%���G�)֪�5�PLY������䉺�k���A ^^]���S�}*����g`��ma��	�2*&@oCu���9������X�\\���u���� �Е�K��������'q۟M��[�� �J鈙{`�؞�|�eP�~�!`�{j&$�B>������ 7��*V�|����^�e�1Z	��d@)�B*�
7�z�ܪΙ9
�Y, ����cb�++1"�{�[U��*���P%��Qi�[���7`4��9���<���F���5���똣}K#C�M��v Ͳ&7j���fc༿�l�?]�="��9Ʃw��pjՔ��Rn�,���:+�=o��OmװҹȶM'�Rb��'�)�IZ#ү�6��;�b�蝦;�؁'Qi�Ln���^�n�x�J � )���X�85А�����~{�:�ħvP�*g��>�p�&q�jz�t��Q�r�54���+�3��tY�@)1;mv��ۑ�9���%%�||��})(*~w{%�*ή�}�\l���͏�V||H�����oSY(H��|��M�=��]���z�v���RfP���ņT*�"�qܷ�oqyݶ4:mU��z#������v��~����H(���[Ι����,�[/����;�a��u�*�w�ށ2GC��M�Ӂ�ZY�SPVfm���Yy|�`$;}�����#퐸�p� ��6��/���K��dr�f=���J��8�d0f�v�Fd�:��ߤ�yw�<��Z*���-��<����F���_)�����q�Cߨ��i�g�c �J�p���?I�,E��xc��Ν�"wHRb)�%�DSL�G(��9�h;��B�>����1��$�xxy?~�u�:���T`���ݥo]�i6!�~[�ef���)2$j6�W�����'?�"�����\�6 �q��:�|�Ց?���	�S���J21��ƒm��JpXR-�;|:|�DH��Q	�+��h2�omo��h~��؊��OY�����wL�%q+�E�լ�WM-Ä�o��ڛڡ�G���.��Mϓ��_6Cٞ%nCY}�ȟ'B'��k�s���I���Cy��٘��ʇ�@k�+\�ͳΝ������
LD�R� ��
IQ�M:�{{b���溿z��^HCD�`�]h��ma9�e�E�Zd"��:����Q;$	�?�LW%�PN����'D/�u�ۦ�nf�AY�-u���\#+���b%)!��m�B�k&�!&�o\�b��g!���屍uSȶ�PJ�ׄ�āS{�jj8�P/eT�����<@w	�Zȵ��T�: ��.�z�s)�w/
��h�4HO@m]��%S.�2�s�UUU4�"bF�>{e=at�y�\��Q��~���q4vpy�>��J3!N�������nJ�&���⾾"�.-�c�Q���,e|$�=Wc/�tH��A� �+z��T�W���F�KMG��8s���Jt����2R�<=	��L�#Þ��؆� ��2�f�j�c~��`�{���ze}�j�Bz�v:n��k�}���s�wvv���p����9�WA%Ij.9�y�jl9K�62;*�^z���r�n��pἽ������IQ�X�����x�`#�[?��~�?�2K�s���d����`���ĶY�È���:۞���i/�6|ꋓ����Tj|������×] i �/)@ġ���z�P ƚY]NB���6�H_߽E^Mg����|oHw~� Bh�?1��p!)r���������&<)(#�g�gO�:��M-��^Cv%��m�U�_K�b_�����`A
%�C�X
yx��d1���uﻎ�F�ZY�ߏ��	ԧP�� j�M� �����v��W��A�<CD�ߐ�nl�w�tnsG6[�d�ʹWJ�i�Dx큁�����+�;l��^k4����������
c��d̫uҹ���#�ӑ��_Eo_��4�4H�NMM��ZLXk��/���ļǅ����eϥ��������ݣ#���i���?���~Ki���c���Q�H�㋀O��廪�~\�Ý���^�� <͸ �X�
$xcz*8�%@y�:a}�433#�y, ��p�"���nx�7��Bw��q��so�{�<?=�$�(f�= T��|�ř��������9�&Y�);?wz��?�#����u	�Ə��y�KHo��H��v���V��v�(֯y+8��lhk��~C�f��R��^>��FrQ6u�GM9����8۽������NTT5ZC���A�n�e�8��#Ԑ������!��x�{4
)}�	���R�!s[�Ĭ��0Y,B�rn���;���:��d�v��!cq=��Ǘ(������	j 	Cɕ�u�xvQH�M ��/]���DJ�+���C��e,���� FӘưj>W���n��6l�����G"���Y�T�lr>��4] 8��$�Т�����n�V!2X}s���8<�F3�&�lu�t�u2��@���}Ȇlk7����Ϭ�HCm����0Ʉ��ev2W�*9*ܳPv�Ug*.1�Ŕ.���5y'Hc�FP�gG&�r�=2ĥvg�R6�{�M�V��1Q}��ʢ��B ���͋�ӓ�l֏�]=-��D�"縋�T1��Pl$���C��[�*ZN��6[b��JrsN��>�M��ٵ���{ N�FxTl,k[;y�t�� U���Ⳣ�-ch�Wy'��LP�+_\��ZӤ�c�.%�ܜee��)Ťs�[��9@�f-�^kK$e�6�U?��G��&%`�������D��!��Ʃ�x&ͪq�D�W8��0c�v��f�r�r�Ѥ��~��v��T	;��&t�������Z�Z�e9�f+�49�u��H4���eZ�6j�5�.������Gpt��
oἏ��zB�[�W#roܞ�&��|NNN>�t�:�����J+�Å���۹�e�멹������)7ph��0�-gʴx�g�F���Z��"Q'B�8S�&�|mNC�v��#lrrR��6B�������N���`Շ+����6�L[��i�D�S:ߩR�_�#�4�j2�^���y���{B�@��'��/�kMz q�1t��	�u��竌f ���/���)5_nÊ#ɡ�_6��I����#"����ɸ���J�lƸ�浇��nI�X������{�%Y����K�d�����g�x�&f����.�v(~�e��4%���,�@vT����x��}]@^\����{r"�*N��aww.c":��|6po��}εu��� ([o�u"'��X}r8K�1��<u����~�:�]�|yd��M��g426��1��L�(�\��é���{����Q֝�Q�S��o����s�ٞYc1���@;5 _)S��WGZ �����W7�ϻNo��9��d�=��l]X�R 9�A�@�+�t*�R6#�s�sh:�%
�v#_��@=�ʓ�<^2HR�=HQbAV!�<�>2�S�s�o+��\���냀tC���1�fl.T�풄�hv`,�Ւ5� ]���?��7K�V�~��κxܷ����8�I�K���	LD�]�h]Q��=�-��=��˽���c�s/��KB��C���g���?4
J��c��"�o9vƂX�%�>�ޜ�'�=>������DKC~��A�a�0H4A����l���l���#=Qc1TGn��%���~cV�U^0�i����o��x&ͼ�{� ғ����t�Jғe;9U2����'��,x���	�`J8�xqmAR���NPKr��ײ���h}�Pbp��\�������*dGe9׫�'.����		}7�_0jXĊ��J��g[_7 ҹ��n5^.�͇u�9|A��X}�h�3�+f|]d�D4�ߙ���'��z��om;1���oH���X+��"����;U A+�u�%�����. �$w��-3�5�'(��=H3���^�R*�����
���f�:k�G���/j��d}ʾ�SA���y�����i ݠ�������#� \^]1{f'��Fw@�*N�w�~�KkZ�]w��p���@���C��C�a&>(_�����>7:�d���ȵ�@��^cK����K���,���;	��Y�W��$x�����9�����3o�F�Ԟ0U3�x
���9��&��k���F�2r��}(x��vJ�I@҂|_7�$�Y8��P�N��;�n�C@�n��L�\��m:�@݃�����&��ӓBH�Jr�7�$��l\\A���n�947�Dȧ��܂ܪ�����
FQ]�fEׯ�C�������IE߅i\�o<��*Q� 8��D��R�Ѷ1X�.�>��s��PbtK�[<�FU����@���.ϋO:��F�R�l�� �|�c��9H
�6��r3I�Q��*x� {����.v�jj��"c �����3�q�B����2h���s�n�#��P�!ЃU�FA��[=����[J\2�|+$�J��9{2*L:���B��O���B��KjC;�zρW���	ߓHזp`�>�!�Ѯ2���X泻W����u����R/�����7IO�ȯ��'ޖw��d��}{���G��8�6@��!TĢ��H$�~��S���sBb���l%�BJ�8rWjK��:�Q��pZE�� ��'��Ԏ���m���o��Q�r���ң(Hq@ۧ���%���C���$À���X]�0F0��D9�y�:p*��1��@�F���hq\`�!P1O��*�椠���Sj?��קp��xR]�/��i
�Bk�1�%����rTPV�����ϟ?)K/�Mn���:�>i��4t�!�wQj��O@���1~k��;��Q���y/�����&;3���gLx�!�P=!@�Q�QY.���ZX>�6��:o�N��AƖguH��M�ߠ��p��CyB�@~����Y�_�&�zr��۸'�;�}q舦��zt
�:�@�&1@�?����w���^�H?�!X�Q�p�'�-�+������p&\ �@|�ME�\Ջ0r��Eh���s5D�l����:VV�����Vip/��t��v7�r��y���	Z��74X�/'}��YW%�@r�
��0+��w_l�Z��O]��7a,��bH�$'p㓬��|�j"ݣ�$�7�̋�:�s���xxx &ym.��$$�rP�Gvm;t�9s�'��U�+�{5yNE��� �Tj��c���Pל�*\�1���� ��]>�<�k�t�yxV��k���_��`�����'�ߗvoۏ�|�@��-B��A(@��y����ls��l)�z׼F�[���&�I'����%S����?�A����fB�cBp�4�zF.0�Ho�]��/;:2GM�� ���2�&&���5�9�ʴ�V]�
a�����O}�R<]x���J/��ȴ���G{4J.���<!��;�{gvr�Y�ͱ��W����A'xs_�����Q��/���p#Ĩb%l��m:V��R���u�e���!<�?�&7��~T!S�Svٟ�z��R|P'����A�>�}��ˏؤ'#J��ʔ�K���]WnE8-����.h阾���2W�E-mF�V��Dè��d�rm[��x3#6�#H�X�P����0U{
S���%�f���)�z\J|�@�F��B�2����1z|\h��9N�R*k.- �!�#��a$2����s Y!�G{��2���t�rs�Wεx!x�uO����l�F�<Y�+Qb�m������N(D��춺+�a�y̲�����9j�f/)M�L���-%#)
��A�,)#��O�G�=e|�]ZQV#xB>�ǟP�Z�1���[��������:s#(3�^:� �����h�Ԏ�;�۲U��-�nD���UZ;_s��ŧ0帻�c���=_w�o���<�����sʘ����Oϙ9�Y�؉����K1ضs�>:%��X������d���5��٧�8]������@��8/���K�r<�����WN��y�����>���q����/u�M�JX����#bG���0"�ow�0#	X���c6����Z���,5���n��O�iF�y�@,��iӉ�V�!���w��$c�k��L�3K��c��t�ي�F66����k���|���}G �T��Q��"�7D"+�"�,6 R����U}?��q�����[��oé�l/�hWY@a�p�݇@�<\w�Y�"ԗ��*6���3���7
�;e�ڮb�m��0�7a�o;5NZ/�^�^���h�/À��(��<�8�~���4\��B�Bz\W�н�n9i_�(T�k:��hk״O:E����t=�~�	����	FZ����iNEh'�V;m�_��j�w�
�P^^�z���|���@�:��v�U��v�]ߥ�+Ъ%��b��	{�����9��<����nM<�}~�=�D�%%����e�0�%V�����Nkr[�G|�Y/۞w�B���7�����&�����(�T��8|OR�9��~UmM,C�U^����ol��mn��
V�n�d���*<�
�%J�h�)}��'f��{�� l���D�a��;�#��%7�~�ngj���vv����`������ͼ6%���*���s,$�v���-���ڸ��`|�=Я���o��]�l+�������>7%~�f�a��R�q)nl�����q-}�ef�����m^Œ_�4HP��	���^v]}b���/�[�-JB�"�{r��r]��c���Gf`<Ht뺅B۬\�C7s�B�AF��U����*Ha�cq���ܚ��'���ˍY������/	��U�vO`����x]s�[ܕ�D��r/��KK�9323�ݵ��H���^ƚtЁ� �K�[�9�G-�az�F(��2�/R8au,��g��>��u��n0��5^��	��h��ֳ�GM:��.G��g�й��,�E�~�����U��lSn	UKE$��I\P�g�e���+�s}x1��U��iで+�L�5g4T�n�G}R�ͤ��Ud*�r�~�߁2�����U.��XZ	�z>���Ru� yG�Ą/��#����ؽ�^tad����gi��[��ۍ�(vߕTOl
ؑb8�����ǣ��O�-�ڕ�_9�OGC\�_tB^�o^��_![g�>cvЊvq�7z�gM��J\��Z�AN�=������-.YK�ZV1�G���;w4<��?�9��i��#�bo��	�°g>i��_�-��w2y����t4�@#�'m����H��s�>�E,Y�S�L��K�J��*�c ��D>3T_��***�
��W8�c`2)޳"�@���n��-�Md�������Y1&��̌������g�͖B��;���n��:M�o&�>�sp(�~��@
�����_�z.y�{ Y�X�	�䠲�њ����FY���FՒ;A��#2�J���Mda����5�w7��5�$000�GGR���:��nή�F�?��Qf@�Q;���OU�����{bƱ'�Y��]�|�V���Ό���,��j4	C��?2��*%"$�;s*�a�)�ؗ�G�>��	��e�C\��R�s�=�RI(P�]N�z˽m��_5����D����:�>/�uf?��{BQ�����E-a<�6��>��?�?��u|�9Z����=a_}���}% ��^��>#�f@���%�1�3�rv���QXQ�,$��fe@^�W1{�>5Hcٹ�BT���P!;p�3 �i\�V��"=��P:�3IT#D\\\_**Ї��)Y��D|k_l~[���


Ԑ�����"H]b���e>gp�"P�d3��mF]S�z���Y�U��gE.kNA��+�v����ZV&Α.I�v�(e���BDDMR<e�� �p```�pi��
��o-�o��Ym-/�V" ��:�����X�'�O�J�F����Eb&+����/A&�����**��31)L��CH��w2x�ɩ����v�#��؎ε!�җ%v$�HI,k]h��Ob��� �s��E��S��=R���ԯ7�R����������\�x7�cE_�^E�߾��������y�F��o���
��I0	��6j *�Ϭ��ef#���ׇM[����p�SL�C�2�u�m��>z���#r��c���T�y��29�nb��+H���A��in柞���G�#�*L�`p�LJ�7?���e���UӉ�1Ϟ��R����]c�BY���,	�f㼺`�dm��Ey\ұ����]�gXpQ��E0fX�!�������Mk�8�ƒ|��L8Q�� v�xд�_�?��fQ�3�m���<���LJ�;�|�1��o �~��5���8/v�z���x\������S��O���L翿��������
b*:;A�xd��Ĵ��nU&����!��w����_���4k�M{&��#}��Cs��x'�p��m�Lyfc�=Yȥ�r��.����[��?Gը����6(��n���9H�$g/Z#YZO���Bߙī~.}�� ��h3i^���i b$�7�kW�.��3~~h�n��R�2��z���1�"wH ���{�¾Y��܀�c�CyfbF��&����-��?~��h�n�AؘB:�58�Ywmu56>�7����8���Ň���hw���e�f�)�]�HX@�x��х�T-�V[̨q{c_=5~y����(�?��,�
�I�þ����ܼ�JG�
\��P�S�(z{&�����,;�h��{;−D(U��=���X��(<�ȳ&}f������ܬ�5#��t/�\ssq)<��)N�����tQ�M�zn����w��Ķ�Y޳��6�T��|��4<'ze!�:2�1��`���4{O�X�= ��}��Tk�c�+��?���[��&DO�W�YD�̽�퍸 �/���Ig����`��:�pu�]�����W�U���Q��Ǯ��4��,d� �	砥�9G��4�x�b�H(h��&���$�^(U���F����y�$I�cPkO��S���s���m8�)�C�^*+1 %L��a�!K��EA2�3E�����p��(��2��y"��	Bp+���-�e�EK^Ș3D��cIR�y ��)��1Kԛ�dŷ׼��*��,\��Y��d�49����E	�.��J��0�����\�`  �7]h8�G�+��W;���	�0Z,�4H]�6[��f-�*�2,��ի�/I���ǆI����$D�έ�c�g�,w�^���Akm%�GrE��׊�U6����ճ�v�t������-++�������x���;������{zz8���*;m�1�<P
�a�]@��l��d����%�|Ez��+p����Zy�r}i�H_C��xK�D�(dX?Wt2(�Ea�P�� �=Cɔ6~wM\+��q@��`n��������w�)�A:߁ȇ���t?#`�}����&���]���<�ô�����Z)W7 ��mF�[yO?D�mEE�QD6��)hi�C)��f,]���;�B�%Bw�y?΃
S��Zl�sێ�@�/K����b�P��I�@U�7f�^�>ex;n�Ȕ�!cS��	4�7�B䇺;pm��Fr��d�ٻ<��3؛_!1Ts�ll��̩B�yZ���5��u/O��ڢ6�*��1��GIRbNyM8/��p����\tLAL����5�~�3�H��ԃY�����z���q�t��)�����+��4�������]���䤖F�o¤K\7�0��43錪��K� ?�B �μ��_�1�?h!�^˶�6��
��.&�����F��Y�ʖ/}o� 	��;��������0��!�()�L׻�߁@t��r��)f��&��ֆMq
�ǻ������so�̂�an(#�������	9)��n��Su�����^k�N��$��'��z�j�S�4u�g\���H��	,�0��HMB���GH9d�j�g�,���ת�3/�1�_�mk�wʼ`�C�TGLC;b����� ��{W��ug��C>��6s���x&۷�Z���ON������"/�1��κn9��%;��5��z|�>%d��XHaI)���6��Yj��������15���Q-@\��J�5X1:x�������L�FAii)����f��~��U�(�9�{��8"%N$;��ѢM:ǽ��9%$�
�3P���UR����_!ߝ"h,�s�4<�d����t����~�����%��%�|��_Q�:��D.���	��:.9v_�_Js��
TF�~�ؠv��L�P�"_D�pjV�0��|H,��Cڜ͎��z�������q���� ?�!�������k��KW8p�ox-W�֦7�{;�8d"G΄�2f��|�k_�Q�毬�o�)�$$\�fnE�ԙ��k�YW���)Z1�k�p�����ي9	�|F\��N�u��*K����ܶ��~�؇��7���h`�	W��ӑ����P�yPq�UFA�->�+C<��u'��ۈG��*V���S2&%��ɚ�NZʆ̉�s�*�����Y�U�L3�����L��_�K���l�0�=��/c�}��˘x���@��ڎ�K��{n/���ᯪ���B6H�'A,�����BA��ߔ�o��r���p���p���śY�,5vΨ��㤘8;;9	�{ �G_Yq?0SH~�t�����L���i�l-�Z��[q@��C�Y9:t�~ӽ�4��М�ן|����ʙ�����/0�u¿����I�J����5$N��p��H A,���A��ɓ6�E�����L�hЦ6��H.��h�ėH�T�arq1ryYhwL�,�"n�R�S�M&с��b8Li��QD��Ks��9�q6��SN�uB˂@��'��5�x�F���6�J,�fc��O1���K$Ss"~0mN��,��5�a4�i�&}��ᦦr.�/Ӿa��i@�g,���yBB#�4[Q(�:�CI>��:�S �G�ӡ$]����F�4�P
�5�蛿�ǉ?|��Jq^���W=�Y�8��"LJ��x���l_�5�2ב�3��z�	!+۱rX�fx����"Q�趸9��[�Z�*�P��ͨx��Ge�PX ���,F�?����3�%R��@º��Y�<#�ka�̴��Vx�V7���;���'��������zV.pA�T��[a�&�5y%�P�la?�pF-V-�����(��	Ϙ�d��e� #Bo=<�:��Gj�����W5tXSH�]m���Ts5�J���}�ރNA���#$b0!���?����g�:ʓ�<=���"7#z�`{K3:ԡ�#�=FS��� 2[5�N�4�.w̅S�q� 0��O��'o�k���:��T�/�9@������5b�n�&@�:��9r��^�:����PPۇ+t��
�y�_�@�:-���m�ZA,�;�5=��+�W)LjB��5&3�X^���w�j�:�l��
�Y-ܝ�����4I��9��-x*+I��B�q���DA��O�?%e�^��v'�a$@v/]�;,�ʯ�J�o�(0�ʃ��5�	��T�����@	ǌcw#��hR���H"W�X,�a����[��Is-�ƊȜ2���Qi�Nv�Ci�W8`�L.V�J�a��	Jvɏ��C޶����f�M�qȫ�,tf��=f��F*�E*Ѩ��������'fgC���[�$}}Eb�.^!�.`E���b�3g�����ˤe$���e��4���S���#�_��"�	[D�NGZ�.�d�Q�H�Y�%�)NNN^bW����뙦���@��H׊s ��.��e��]��!]�j�������OF�Rz��i��$���ϭx����J?�VD���Q�=���W��%� �!��!��1��-��())�t��]A&��IW��3�K�:(<�R���Q��_�_�Uv�~� ��d���Qv{��)N,�{��3Ƶ�u�Z�a���'�k�Zr�z�x+�k����?�o{Q�����Pt03BܘR^���y��cJ�i���H��s��� ?�=�oo,	�aM�oZ��K�v@X��(���e�ۊ;����tk렐Z�9x��C&oVH��#�2�Uيc{Ӌd�*�	��o��|ᠣ�z1�Z 3���>��#Fra*^WK�?+���w���� �)�S4p�vZ�۔q�᚞GԒ��Gܿ�����_�P����l�x-���=Q��	���e��Q��B� (��B�K4Ѫ���'�3��-ݳ����r��(i|��,�|f¨����������B!}���&��!��ϴ�.���	h�3�W���d�d�d��d��@Sww%���CI6�`?Ml�	�K��2�ߛ0���Ɋ�Y�X��.T��)/���eP��#<��1��2��!�W �Z�t��÷T�z��%g��bZkE�o$>7��������)_�Ǒ�+�O;�1^�tZ���[�
��N1�9U~
�B�0>�<�7Wd �'n4 l������@�4Ux�l�p>���x�H�������P�%���%|�,�5 ��Wc��+*W��>�����bF�>����}�rcK�׭w9Z0{�����H&y�7�-�V�p��pc��m�x8�jy\ޝ��w�d8��L.�s,Ч�~�@h^��4lϕ�a'LP�ճ�}sF��q�5��"�,��c6YR�z��fnja�r%=(3l��B�n�9JVe�q�)�J���m��C�ۦD���쌏��'Y����^ /���u����f]Q��-�+��1J� A��x���?财���1��d��rI���_� �ʹ\��\c��&��8䌬w�G���~���WQ�r������ ��Y-�2 >·��U�*%?���X���P�a��(�/N���&Z��Ac���Y��PEU�R���Oo��T�µ{w*$+�J~� nv�F��Ψ�+D�`�A�	�G�n�)�UQ�ht~˅9�䀋
�t��I���1K՚`�!�`'� Q$���Ϟ�#����<s�[`c�'�Op�&i�	bø��(��(~�VS�X�O��b"�0�%M�K^��ʴ��S��U�>a^_g[В�/��6��D�- ��x�l93�����PA�9l�+)>��z���`����g����[�k
�~օ��S�Cb_�����7"YPF���kcb�h��0[<P�嬉�n'��8����;�/d�c����b�z�NP��ޅ-)�r	��I0��xi����xX��r�s��>m�����ε�$�DD��"�E-J�����;�Q��D�]�6J�ha�т轎6�#������>����{���k���Ȅ{�g5�SÚK|����y�'�no/�遳&J@��*_�:���1�9�v!$_@�����!�J�d@LQ֋�w���� U�i(��r�lx�M��U��p����)�%d��V>���K� �O�;>8�TC��b��\��$��9�������7xy�c��"Q��d5��s��~�A��-N��LN�d �IR���@�NS�'��������ׅ��l���Y_� �?lB��yw�^�2'*5�(�Ց��-����ng~�`��`�p �T�� D�-�,a��"�Rs̉�IV>h��6����*�����!w�[���bx�a�����}r�{z8I�$����
 Ʒ�Va����o�����ϯ�k�䳉ט.f5��9���, !���A ��!�	Oʇ��ĸ;�x�C�h�z	m�]��5܅�G$�� �=ȁ`K�Gu$^6���S�R�Y�E�Y����Kc�����I�t5���L7"�s/�W4r�?P��3�`�qO�f �;�C�?����e�P qH�>ݤ:%���ѷJ>q-}.}�M�j&��r��[�+�-�y1��Q���O/r����L,�|?���
U�;R����q�Μ={0(i��t`t���ߐS&���&���ۍs�oO~�"�� 
A"̀��w������\^G<K�y!�\6� ���&���>8I�~L 兵"�XU�h3A��<��@U����ZV���H0\6��Fdʛ�Sz���񄫣ף�S��9'2�W�^Ú�r�ԥ��u5K_��Z&,�-��������M?�}���?m�S���Y�<%�9����vRki�g�Yw��|Ի��%'!Clxn��~�m0�A
Plp���%�˰}��D�
��oV�Q��H��ER��Ҵu��
��K����{�
�r���%$�]ox� ��\$C�P���1�,�,�R�q��@#h����O�237D�"k?> n�9�x�PXwT��¥��%�����I����~�[�3�q��6%1p~4�[��":1H�K�cL�|,5D&��T8��^G�*�ǟ߈�l���]~.�b��p d��/��w��E���2�|_e�Ȝ�V\�d�`�����g��'0	��Ck
se�j���7���,ֿ�o'*F��W�P�WHѱ̑�޸殭f��N�.�+���H�>��h�s%F�u�	��_�d��+H��?A��^ה! rZ��,�2�(�~��ǿ�3cus��o�T�Ix{��$��r���^+����p��#����呡�1J:��;�\\�H[�{��ب�z��
�ai���%<K|x����7D�㼚���Yo���#�)��U��:�>�ר�򏁐�zd5DV�#�)s��}3���+b�~Ne�35��)�������v��zg����Y��1]�k�{�)���mB5f~|���&��T���#IL�X�mH��l��OV�8bCD��3;����Gt���<�T}���{���yg{�Ckts�~��P�%o��ǎPV����	�%xG�s��NAI�i�e_R��!��4�)Y,v~<k!,��1��ah�ښ��a��ge��������)� ��d�~T �H[����WĹ�SƯ
 b,k���BDpӕh��.鋵�Zkx�C�ޚ`r!L��m����q��ǶFr��^"D[�⌸2x�%WnH~l������Y��{�\��o�J����G�ZJ��\�gɅ<~������UU�h8+.T����}�H(�� "�$�L�n������r�9��+Sׅ�`��Ef)��׭-������>%do��@�x�Fm�s�������/��vnY}�	G�R��pi�r䘂�s��{��g�����?�7�j@�<l�ueN��\w
�������uV���m��a��k�����D�K���&�i�s:�mp�m�A$�T#h����Џ�7���À/��p�&V(U�2� =F|o< uH!�IQ�����k�W�xs����A����=dD>^�,���`�P)J,�}�I�^Gۈ%��	(~Sɞ��0ᴑQCԝƀ8�p�/�tNǖ�����[Kx�:��9�Β�+���u^Ѫ��El�Lq�A��w��`��<�
�,U�8%T�c�8����ӘG�+����%�jM�L�;���t�6���3�---M�U;�u��EyMO9@��v��i�L���������,U臢c�	yI�1�T�����¼��l� R%|�4�4��һ�	R�,|��ܼ�H48��a�����DȬ��vi&���z!�_*R��~�:��H�5�I���0�aJ�	�rΩ�n����h�����y���u�\�Z�D%0�6د�US*0H:�!���4�fn�Cv�����'<�=�L�r̀6V1��uYh�����X�� ґl�Rm��B)�l���q��<���įN̨�V�����|Gl�黀zp=w�u��n��+[�^UO�uIV�U�qR��o+J��O�P��e��y��c�y�l��τ[�Ʋ a��Cϭ�=��e��z.�����ZN��GN�u�o��Nd�ʋ�Su��U\�����U���� ��^ ��ஆff�<�� ��K�UB�/bw5Oϫ�u�$KA�g	�w�TR��`6a�+}���V9r_���
��S$x�;�����ؼ8���8Ċf���$�)7DH�m������.Y6�񽧱LŖ�{�����Q�zW�Uz���0��I���ҹ����i��n�'�DT��c>GIj֓�W��'@J�k�iĉLjp�(���yo���C~�/��H)qh�bp˲���q����L�	Li��U�n�_a��F@��M$���9�"x��S�|o���iL8/���Oۉ�r&�t�L{�)ӕS�m?a�'̃��-�𰗧�Bh2A;R���k0���:����VN��g�U��B�R�+7l����V8����x�p��lf�h?�o�Xv}��B��M,Տ6h�$Wg�}+W�P�~��yˉ��vPK��G��[�����K��X�����Qp�����g����H�޵�#��a+gF�����X��jݙ�C8���ӒZ%Ͷ��;/���U�j6��9$Y�4،<xv��;S�0}�iW7Z�A�𓄈���?�KZ���7����kң��B6���z ��$S�xE�U!�3��w�8����<»l�	{��5g~���[%�����ؠt�e��G�b��&Y�+�Q	/6q���66�7v^-m��V�ӿp����n�x$��ѕ0�ל*�HT���g>�I`J$E�����un�x\�n�BK����cޮ��PH�����Z�f�v�.���=�UP��'bA�48p;?�I<5�-Nт�ͷ���j��������$kg�?�Yo
�yn�W8�g�l<�#�k�K]
jrn�)�����������bq,X*,D���ZYi���Pz�4(6��]��I
����b.���{Q���E�*��]�����+��{�/4ǡ,��>'+6)�N�S6�y,�}a܎8�v��b������ /{�8�p��$4��w�*�g�i�]�f!u�d=qi��on��wMI垝�"9���$�~vg��[�G�m3�k�#�$H��]�=>O�T�^���8r��j�T�&z�zϫa�cz��:�ƚжݧ0�9�!E�VǢ�"�Pwا�_%�KI�#���X�ٿ����r4��hߑp��5|�3(s�N�����e���[��+��dL�:�3�\�?E�����	,�J�D�Ӡ@�QK�x����WH�^x�6jإj����G�v�����E�b8N�OX�3�(�q��2��D�K_��pvRjE�d�jQ{_T�74�E�k?|�ΒG ��7��ݵ����DG��I���H�S>�+0��R$�D�����d��gg�j�ƊUh�S1��<�z +�&�����D�=�֢0�_������o��U?ܚ�D�S-���L����d�` >���/�Y�abM��p���C��c������x*}#B�~���Ձ'���\�+(t����5��������P�S#���3��(��
j�Z�D�9V������ޑx)s8m�������
�������`�7�Ӣ:�b�۲�[��{#[�i߮,i�iʬ�^_�%Я7�3 ��!��B��UoYU3�*���,�y;�Ǉ���k?��~~����{r����	��w;K�vC�����fp��Ș��E�¥�$X��)h>vb����A��E�l�ES0E�7X��˹�O#�D�����I_zH�I�7�R��MS�y����yv����B��v4-0"IZ�5{���4z��2>DN�ϯ��O�z�f�G�~�=�:>�:�F{�^}|D�sr��w�#W��)n0��Z1�E�}��@L&��4nc^7����y�<�Ȧ{��B� !�(F��H���Z��"�K�9��.7ݽx4Sg��\�`N�ϵ ������ՄƁ~g���C/��WS �X�_+ڶ���%&��ү,t�7��p��%� ��Z
�ri�~�|B*"��rP�Rq��R4j#�1f{w��W��J��~5f]C��k��r.~�3��2��z�Z��?����3�3�m�.��Ȱ���C����,T�o�#y�2��@��Iʺ�,����j�Ӡ�g(*��l�D&/<F���H�e����|(��3�;�{�gY����]���n����{v�T��~��k��հ�!�!��t�(3vA�;�>��H�s�=�q�2��a��Ej%�j�ޞ/ J�����{H�5q�r����;��X����d^�霷?�e�}	T��x펬LtZ+%�i#���0�D+ekN�e!/���EL�n��,^���4H�'�J������F�����M`��yw�Κh)tG4p����(+#*��E��J����E֭*��b"m�Fѹ����h�JzI���	4mԝ����� �>>�t��i�T�&��*��KbS`�r~����v��p�⅟kv�Y$�m��#�m�ݟlm������9{~�����R�����1ϻ�;-�̓�	�ͻ��F�,_�K��_��;�fm_�.�f�|?0���T����(/'�d��|��3� �~/,�k^���	K�����}\`~ZS\�Z�~���K�iu�~�ӏ)�%#}س�` c��@*�0�K۳�5Y��2�Kj��0th������$QV+uUuW�ũ6��)���1�r�}·~�뇤�/z�'�c�	s/~wȔ�*!@6���C��n5���O3���y�8�ծy�ó���X^^nL�
HqV�b�F@��x�jKK�!s	��'�������g�����6q3����O�|�/�d�G�ttt���(���ٍMf�&0ڣj5�j��d��ϹvO�{�i�C����Med,e���©II��Un�=���]2���nԽ�p��l��g�/Y17IF&��IePx�g QW&�;�����'�a� K�>�F/g���@��~<�Ho�?l f���G|+�$66��U�G�Z��
�9�e/�vo�ud�61�_W�<�ݭ]Q�눿PTzz��B�F��IH��P�r�Su�����t��?�F�Ww�t�U0��SB��tl�gW��+�IC���qE˹�LX5@R��A!j��{B�"ڥ{�n!$��%~Y�F!$�~��x���-mp9w��s����8��@;pQB���|S<����G&��e��avE�;�iJ�gĺ`�H��W�۳�r��ץ���I��}���ˏ	�i�� v��`YX�B_�4,���,Vg	7	W'kMp��#`�<|wiip+'ArX`_eD�ش�W�vM)G�+;J0O�}�.�`��|vDr�U6�����(Fmf�ͩi@��#�vK5{��*n܀ԑQB�L�pwo,�E��1G�f,9�[�}���)�M��4oɿ�.��O��s�w�C��K�ل�"��f��$&�s�{��*L�e.:�𘅼��7u���BS����U�Z�8x�4�Bmv�0��;ڀ���#�6�����ￆf/���7� �x�[  �t-o@�cq���U�q�d�8��]���< @u����k��n�$�_ Üs�Û��r�������+攝_���eb�k"�/�MP_.��]#������H匓��S2�����}I[[�{������T���`/��H+0ᵅ���;�S�E&;�J�5��U!�9%A3lh Z����:-&1[�T����[hH�ܜ(��^� ���y3d'ʔY���N��=�	B%n��(��!�Z9��t�m��j�$|)�/�L�7�B��źz����=%W$$����2�@�>�M$�Rd���Y$�rJu�x堖��+#�49��Fj�z��y�l��= X)���^��"���OY��%�SpBm^�o�j�������+�е��\^���E���t��W�8�fu%��=�Ԉ��S�l��l�Ŏu��2�K�%�	<y�|��I���?�q���RVh�Ӻ�+��w��2�dHh��E������\*I���S�ܒ��C�ڞv`K��t�H�H��A�E+�Zos��������S�<[����nW��t��Zp� �z}���}Q,�(ϗ ֩ۄ���(�3R�_�eOn�4�?�TQ愠�_N"x�L�Hu��J9��YH*ć}S�dp�����3�O6� ��`�p�h`p]BjY�P���t�O��xI��I��'����y���]��E�:��VNo7�2�%=qu���.��B������	a(��W�#�̊��@�Q�����(�e9ۡ�yQ��h'�@�\�`ޝ����s&ƚ�@��W7t�!��ק�r�A���]�%�nPJ���S���hK4���1�/��y3X��,�I[����Vcq�mq�Qc�ת���NVv����J�S�~�-��H���T�a�A�a�^��j̜D��Gb�\�+�����%3Ͷ˫�y����RfN�:7��#֤��9'���x���ɣ]������̸�|OiCO�,�y�h7Ck����#s��sr�$K�]~�:�_��~}��� �Rvf���g������i��l����v׹��Z�Oq��+�v޾OW%Ѽ�z���W���wL��a9�Zws�Y��W�����K���f���#Q��#��+o> c�S��)r�ۮN��pb��h&It��$���ؿ"��=:jkBK�K\�[g��z��^�&�mP�K�H�sB�d&v�<��m�v8��t(@���'S�8���L ���:��*���H�Tڒ��+-�9qp�͹�V��$=Z�I�,��|�<���t Q���p�_��J���ěK�6B� �EE�>�lki�#��kfp�V?������ߴ�)��_��u�s|*!�uj p�#���/��B�	�g��)��n�P��ig�3������������R��@'A�FGt,�@T�@Wi�	D�\�E8���hF|���x�������g�s
��F�s��ue�j�.�5ִ֞��܃��&�V����/ �J_��6�)⟬��\}G�?���8k�!���)O�@��[W�RJH����m`E����ޠL�ߊ-��	��uR�ɜ�¢����3��ka�\NB�ݿ9�ɞv[�!�D� �{�R��ǻ>�5Q�.��s���|����!�<��;�_�#��l�9���� x�	��zmd�ڨ�ċ��+|(��c�)�12��"ӗ ���%���uL4.�9@�@�>�=�O��M;�d��V�zz��k��z6��=��"���Sj�O�����Y���c;�	��J�R���OLpМȈ�- �o����5��=xo���cN�2��{��"�ӱ�p�ٚ����|y��7u��w�){S�SHvx�L�<����4I�h��)����U'�ojH�kd�?*�Y}�� �h�i�ƿ�{g�ÅM<���;�=�8� 5�!^��}�a�$L����': �%�&�S����f�u���9��C�9G/r��{H	S��^���쑩+M���Ja�/�^�yr��nOXܫ�4\�H\��ϯ�Yð�)�<���L��O��<�~���!��?�h��^D�zs����N���kt�}�9,O�";�dL��2�#jt�܋�;jXd�a!�|����sCD���M�*A��N�}�|�`���_/�"a�»�e�0����v�Bc��Tc����M$�g������WA2�ą��/�q	��)L]�P�p�J)
�e�y�^�g�^�?����ZY�f�,��i��������܆��zٳe%��������_�� �M�;)O�a��1G<�f��>I"� Eל܂��ã�g��Y�j/�S�wW�u�7�t�H����ιlT�-n8J)�?|]��}T�}/�ѥҸ�Fä��¸a"�0�˶)��9rɹ-����<>�~)�3�K��礑T\S�+�����]��"�(v�P��^#iJ"�$"30GK~2k;�5]&	����*Yu���^F�����d^T���|��H�ۧV��=oO��Q��XI`)�k:��V�G����Y6�.�Pe`�Zd�ZId�ꘅI���U���8�_RR�1"�;N����!��b�nI�{��x�=�L��������0{ִ�ɧ'=�������2V�,���?,]��0����\9�Fam��q�?ZfnP��c��CT�qY�5Zߤ=}�7�q\?n<��A/=+2��x԰^ �������}b�Lf�U���*�Bv�L);�Z�Y�5�ji�p;^�	,��N������(��C"��z9�B%z�mu���,,��\���q�>�3WqU��2�������j~2�YLQO�n�L�̆����"J����J�\6�AB85Mq:σ6Mc�J��+˜w������5��TU��،����!�������m���gfh��[D5��@N�~�1�#�ןD��o���Dw!Bs%d�s,a+�����h��@	��Eœ(���r�R�7�>�T���#��:�A*t��fr�Q�*��ścFUa�͹��)��vm���!f��̥=�ʽ�Yy�
"��\'`��NI";��~�e����v�c�0���#���Пw�~����8��,- /u�$]����؈�&�I)N�1�̪vЭ�U\ Qҗ3�(=�hկ��(d�t	���o�S5�z)�r���R�R"D=[�ۭ˽�^���3�4	I4�MÔ��y����W'���^.hfg��;���s�����k�y;�z�b�/<���'_�
 X$��wL��\d�W�y� ܤ�C�A<�^�Ɵ�s�]U�@�N/��s��5&�D���Q�J�Ә�.ȑ��:{^~������F� DeM��n-�9���r�����o%`����Y��I�9�w�|��5-�$�**�E�4?U��ib-B�����o2��-�e���<8��z�� ���7���d���K���&�Ԃ'c��b�bF�A�jA�\�M���5j�q�1=��K阨F/S��y֎Sh٠Ҫ���xǨ��Ev���f��r#���&"������i�YQD����o��W4����L��,�#�(�־)|���&!yR��9�z��x��n���co��Q��sEc�I����Nc��8N3�������)����j�n���R��8WcE��#\s����b̬}�e�b��v�Nz�.V�91m�� �qֻ�r�����WZ�<?ڲ+.��E�FbC���Q��JC���۫/�V?>+�����z���ʶ�&1���nfNm_֜����-�԰�sLm�M�SL녚�if8�vFUŵ���k�k~{*�b֖���E����� LJ.Nz*0Pf\^&�����t��ɖ�;=�M���Դc�'�8����5���YF��f�~s[���O����;'�7�53fǌD���zy��=I��ζ(��F�e�Ȏ�=��w�E_1��K���l�>`3�c��'?���1�ǯ��(�ְu6��A#��K�o'�f0aP�3�� ���f곁����0mH}h|{S��A��ݒ�[�9/�����P��G�Pr�����+�/O�o���E�{�!D��������q�
�~-M��s]p��c�N��_��9��8�������g�^-��}3��;X��˷[!
�7_nEas����]d_cs�8�-[�Q/׬����i�
�Pފ
~�,�Ҧ��iD4�4C/b�O~��R����L���I�^���e85���|�QCm���k�������,�k��J���]@.Cx6� ��72��Wrɽi���=4�m�������37�r\��4��dlf*4f�i_$�F0��VO��N��pY�m�F��H���e��*�)&�E���ٗ/��o,G�M9�T(|��YR/�5��O.J�eg�Qy��=��`�"�L*��v�[��WW�F��)}�����#��tJ��.�5f���"����	����K^�)�ń�Y�e�E[����a�vJ�4_���~]�h����"�>ן�sJ�X���.�^����s~&�b%�;
6�I c��<������%�nS.u&@�e�z����P���p�H*�45(�'���=��KґU/oU���}+ KʮpF�7�����Y����.rܦ�%�E���gL?#(Z��7�����=�6w����ȝ�\y�3D���7�~)��9z�6�^���S�Y��ձ*0#x��.w���F������Nl6�w��|�����Gis���3K��$���J�W��us�x!��L����F�f��,WGz�J{3�?�������?��6�D�%�� ��v�n��	��d,�X�~5L��Tvz=5��t7�����TE��nm/�x�vc���y��l����5?���:=b�F״��5�X*R�k�9q:\�]j�q�U���5]����T-�&<�r��ާ�!�4.IH 3|Q���\�.���]�]�#��Lc����� '����\ը�3#\�����^�P���&ڭ(A��5�/�I��jz���w{ZI�u��ȉw��I��5j�W�l��^���3 �ȑ3ӈx��:g����G���&����/�وE��D��: �:�R��M�e�FR�_�Q�7��\�����zp�H9��C�ҥ�I(-y��kg��Y3�C$�de���IL���'�C�� Z�_�N��&���XH�s�D��xD��z���a�$;��Y��������ҽ�5���䏻�Q�l��PhZͷ�iu�����Rì϶i �|�NW�T"1>����ƾS��%�#j+�Qkd��U�`�ข��t�۪��('�W����̰Im�ġ�`�U��J-��D>�l��%+��O��8zE��u����E���`l#�>�6W����fTȣ'���ʔ=�N�'Չ�� Sm�sf��]t��b��\a����T�#�2�{��Ib��)D�JZRȚh*�z�a7�BWf�x	��
+�z���r�}�A�gN��)zѺ��f�ڴ�`�FD�?V��[�\�a8\���g(��yS��--�h��26rr�������(��������Ym�ѳ*e�dv��h[��I{ɨ������\	/rŸ�z��u��'^��t���J��4,ٿx��5W�6A�:��&�*�`�[Q��4%��ڿD״{�[MT���"t�,�*�+b���A��jWP�ӕ5�!��>�H�J{�~
S�h�3Y�.F�$5T�57ؿ�gD�˭��F�5���Z�tu̎�=��$���j��E�CL�N���ᘰt��.�F0�f�g�5��>f�c���Z2;��*г�Xu�\��o[�7�q�Q�6c�œ.����K�]��_�]
�;6�Y��,j�ڕ�]���=�@��6z� �v��k�x�����3�o��nV���e�k�w�l�B�N�F(`��Ŕ�j55%̗L��<ཹ#�ͥ��H"���;ﲬ79ӯn#�J��4<g����ɰ�,�z&ŝ�-���U����Tz�&���3�x~ś�����)z�_�HC�5W����OEO�^*�z���X>��*%���Uva!⺿$��2�b )���"l0�e%��̻���7c�F�/���:{y��O��gE��>�|"��6-��L:)=��뻁^Wv�{���%+�o_���{���!5mb��h��l��bK�9��	3|�el�ky�Z��b�$BV2o	�[y��jD�(��ѻME���W?���k������˻ޛQ���D�FŠj�߱��w�/�w�0)��i�gP����=	�tK�iιH[�M$�JP%6�a����|�K�sK�\�A������H��AԬ�V�ط��O� �-?;���R��5b�ܣ�/(����T6�)ϟ�=Ғ'j�*�s��zM-�*\�?�-:�k[�{��j������3>����4X�^q5�7z��:�l���T+��3����d2\��5�B&�jW[|�Kz+\{smez�2��$��X7��KZ(�����/v[���h��l��q-��k����}�E��������`f�`N��A����\�ppWRe+HM"AC�΋e"��@Frv7w����n��f�?E��Md��3�^��^|�n��:��=���=�]�2J\Z�P2���~q ����Y�׽T�sƪD�f�!����HR�D�URۋ3BZM�4�u��c�mJ��������r.�34�)���[R�~���(ql�2 \�jGӬ�85������;kV�Fg�wJ�߷��G�f��:��^YU����i��k��tB��5֨%`ֺ(N�?�.߶v��/���-;��rev=�jp�ތK}<5�×7Q�8(%�um���[1��=�E�1E��O��_β�,~�?�!(��
��O��eS����^V}��l�-Ϥ���Q\�+&���tGj~�xn�g�� o��̟�ǓsGL�ڰ�0m���_t�&�K���,��A�gxw����N��+V�/fVx����Un�ēY��-[tDzv=�{ Y�W��}��Fbɯ-�5��I��<ǧ�"����e�����R����7�?��7�{c�E#��K�$���D�{˷�G>2�6�C�*�ij�p�-�]��Xad�C��c�?$QGY�(s<�����ˈO�'�d���X����q�U�����S|D�����8�mI:cQY��̼�BM��ب��o�g_Ҭ����-}pۛ�+���|p���*37�.�:�Ƈ���$8ު8�B��X��9�>���|�t�#*�s'�m���ճ%�Y�lr�� Ɯ��3{C�O���֩F������6�4hح{\uHW5�=R�i�����m���g%m$��~�R��s���C���~Q���
�4��n�R�G����L�	*_�."N�M-��V�s����p�U�	��;�b�J�xp
�ZUe�j�}f�/wN?��5���#+�:j�rx~�=��YU��_:$Y�)�8��*�£�@X�����1I�*>���<�w[-�jn&N|a�s�I?M�_��Y/�d�j��3SX64u�����!�燜}eM���^�U��qB&���8�x��V�����3,�Դ͉�M	b���%���xGe���^��ON�MiZͭkb�$�q4�\yFs
��N/�du��� �
8��M�L�q8�X�����zH��3���R��z��e7M�Q��3�Zj����׍���Q�@Rb#���~��ٓ��[[�OZE�³��}OϞ���G.D��kZ�<(���"ݐ,f���4 ��b3I��Em��x��2��I�D��U?m��Y<����x�nizp����*��ob6'h�'��^��I�I寊�i��=�qXX�ĠA;�U�e�\6HL�+������--ĥh��gL�^P§�fc$�S�6V!��?���(�<T���OYz	��Ϡ���t ��j,�����	]����y�)�3T���f��dJ�Ta��vH��GQK��Jn]��FL���".��(�;���׃�y��j���n4Fh�]�_Ӳ�����x����Z�ɪ�^�rv�����`:;v�q�||���˲�H�ll�<��Hnï��]7���͚9_٫P_�89���yZc��M��gԡ�l�>����B��:I��݉�'f�7W{��M��bʿ�L�ge4�G`O+߿�q�Q �����r����/o��"_p�"�&���&�4�S�>k�*��ϔ��MC���5�N0	��Y��Ь[����O�3J,�K6�n��;�������5��DT ������=S��d���p�B�Q�c�S�_��G�ElA�|���b'��e���M���'5zΉ	�&M���ZG�IG����,�ɟ����Z�G"�b~���w�)�,XO���5p���X`�%7�R����+'��VY�P��%���cSCַ'Z�8�l�;�g���!�5.�Va���Qm��<Y��<��،>C��}vA��CC{x��*� �e�� l����������Z�ʆ�	fW��(��}jEE�ZT\;GN���ݻl�
��맷� ��G�����,F1��`V��
s3�� ����s&�F��^<W��&S�$M�dw�?y����������oZ�5��n� H<�L�����G-�l�<�zU��N�ȟϝ�}�ܿ
N�h�8��� �#�K(�^�����N��Ls��D#������8���iN4�$n8E#���R���Y��Uř���U_�4�q>��_ZJ��H�r��J��i圭��iD�S͑�5FJ/֩�+%�D�O�d{�{Nώi�9&E�F�E��Rc�xn�
;1cc�	�m�i<,ad?�h@�	��r���S���Q�}��ȟ�;�����X���3/]�RVFƲ�&��^�gŶ�iw&��0ă�G�-��z��Yۭ���\�SqW�{�߄����G��L�j-�l���UL���>���N�%X\��`��;ZyF��ŌV�:�y���q��pW�?�x��u��h��`��Q.�?�����	r�`{D�^vf����*�E�Y�k7��#�!��.kˀp{����ʧL�~m���,$����ZW$�9�h(�>&N��;��6^U%٣�N���%���-�~�u�Y���$�=���� ��"�����`�'�G�C���>���f.
S��N�x��$b�(�޵�ļ��fMڣ}C�=9}:�v,�O�����ƃGO���̠�)�#�ç�f+J*�b��F�"uJԮ_	}��nj�uV#���]%�.E���@�53X�9�Z�xi����n�@�ѱ[���Qc76��9��*�@��*]\�'84�r`�K��Ց]v�~�lA|ư�־˜Ub�
E(ILnN�_s�����Ƣ����Pm��D5h�E��ޮ�V��i���M�Y���jɇ�zi�<X�w���f?����z����vc�anf�^< h6��ϰ|_�V��3�k�r�(Y�ҋ�J W��?���Eg�O���(a��
dH�#_S��
fý�"ECbHՁN�:��AVL��L#�v��p�Xw�t���֚̊b+ܣ=�31�\�����KϮ�M"�|'�h�g����Ivw�0qԩ%��G}(Z�6#�:��-�q��y0�0��O��_���{~�_��F5�6� �m�^��+Z����3\��lO�� ^��g�t�\��j�dİ��b{�N� �QB&Q�ܿ�I��lS�IP��y��	���^G�����k��D�=v]o�-�c��G[L�ݨ�A����Eb�Sv��؜�GE6���½�����y�;;g;� 4�wE�z�Xy-1-�Eu4�~(�Q��`zl�'-�
X���4��`+�)����<�+�H&�i��4�x�����Q���d^���va�Ƣ^���5ܨq��H#O�)��������#�uPb�xH}h��"g�w��H��Ѡx+�)m�� ��y���5$�l���?~y���frdDo���2^Ջ*3D�S�0 �k0����KK�'? {��Ta���"�Ǻ�"��8��ou�h�!X���+P��O@���&�[�}�;{_S\lD�l>:_��
�3>Ϳ�|r��"�8�le�1{j#0I� �4�k���M�����v ��º,�.�9j���նf;5�`���d�l �2��w����K��mYO������/T>�!�"#���Z�����I
���O^?R��;Rq	��z���mr���7[�ۀ%��?��ߺ�0�V�b��9��6�J#��pZv6�G?����C�`�3ZrPAٻ��I��$Z�#M"<w�-��f(]�����C��0!z�n^�Y��gg�Tc�h�#��E'�������Bn#���I���x4^�(��Nڻ�z[�h��^C�Wo�$X
�����T�}Yv���*t]ݽM����_J��.9*����������eVf�2NY �/<���p�}׷j9��3CӐ�N��9�ɻ�,�0����iX���O�F�ڿ����)��>팆�~f_ 	dSn�:ܪd`vXf�x�%�\!�>�B"�0�����A�R����;1�H�Q�k���cTORB�z��̷L��^nv�ަx>��5'�0u�Ā��lBW�,�
����<�m&�:Q�`��M��g��u힧L:5X=v���ƯN���a���lA���x�w@ߞ�9��:��A�"	��r�X�S�Y1ZaU��zq+4��6(��݋������fA�\�3�Y��.�ftl4��MGpQ>��>h��:�ԘV�k_���׾��C���ON��)�hEʚ]�e���e0�!���,-�P��c��+2�c����c섌e��۩��\����s]���]�羟�r��L&`NZa,���6�յ�?��N���b�����8B{�����(�}�����N�E��uog]�Vd�����%��>ĭwBw_�G���އ��UT��h�Wu���M��D�1��Mj�V���Oy��sێ�3���,�^e33�l�IT��I�|�����/<Q�N}\FOr^ttc�&�������w�Un�G%�%M�m���ѧO����+1�O��"�w񽮮�K���a��U-�+�k�����$�Z.�tT���+�ZAs�`���G1��l9KӰ�hc�W����*���>��b{��2Bi�4|��!�]�"�°���f���Õ��Ϗ��j�wP���e}㏞�P���l~���Ş�#NFM��|�zLٙ=p�Y!]��k'K���ɓ;�[��N�1{u��-������ez�ͷ���\�B�ڍw���P�>	:���n&�$�e���ЖRr�=�A� ]��?�8@+��nc�)E �{F�6�z�8�s��G7�jFt���6>�>�ؓL1Kϒ���:�aq$��������u4��e}3g����Hr�sk
H,mV��!�8)Z:���������,G�/�(Nޫ�44�3����A_�>X�o��}�����?��?{��Y��K�����Ԁ/>�rq2�@�X��s��L*�NK�)Ա{�h�^��1A�_�Aίu��+Eߝ��ɨ$�6��}��JJ�	C}�)�lS��NGEv�=٭������Ab�����H��������9Z�W���h�׮�w��S�ڟ ���RJ�5�/s��k���a�~�s�qYD@��E~���&�F���9�ۋ�-qZ��������//o4���<�ZtQ&'u�Äg{�!�lo��&X�)�LC��JR�t�;��Kn�˫���|7\�
.�`��KU����U�6
N��)���S�H<��49�*��e!�L0�_������z̾6|p�;�
S��=��I_�.���?~�]a4Nܸ(��Q�1zS=�WW���C'��"C�eS�c�F��x���m�Ff7�G�=ğ��4	�h��X��<w��w��E���kȋ���E�;��!�u�w�Q� `\�:چ뱇wo?���UY�P:�jZ`BY���O��qv�Ô�<z�#6�hY�
�ש�D�E�{�΅�0�'��ݴ�m���(��d�FT5r��+`ۿFTs�ΘY�w),r��N��tr�e`<v������@��gܯ��q�E[sJn�㈮��v���-�����=K�fcW�R��/8���^�����HE˳LLPӫ��T�F�)���
�i���%�ǈ�~J��s'�${��\�q��g�L��8�3oD��z�Z��:�Շ�o�T��"Ն�!��0�|`�x)KMIO�0��9���T1*�A?���6��hqH���s��۱�=2c��w^�t&6��⡥(�6=p����7,eufDuT5���!�F�(��������<�U�����v���&u�'���]�MC3���m��%u�-kNɌ�P���!(\=[ÅKa�����F�Y�Kg��k�J�	���.ƏE~�^�1��XS�}7�������Q6��v$Tݏ�M�#�R�����9"��G�=��3n3n����$Xd�j���j�P���/��m��Z�lы��Jǿ�|���Cg�l�z؎���?@�Է���m��y�v��\�G�[�G�}!Sz�BI�ЄL�7��#RVIԽ"�7�k�}�Y�E����f�/�?=�Շd�9��a�D�F�|T��������>��Ј�Y�5(�ittޫ�l4X���"������AO,�PVɥ��da�[^D�{,Ƣ���dW ��0��Qswxҧr3��@VYI(�gs�{T��6, ����X�ߐ��ho�	�/$���B�D�?�oįq,
k�Z�?��7��&z�E�1��۸x�*��3�wtG�����;�S�J������x�c�<[ҥ9�	�i#��<�ц�����`V�q�sU G��0�H��֖A����J�:��C�@�5����Y#Ӳ��Z,�p�-��I��;�"m���$v��2<d�7�/�>U��b{��]]ɱ������hլ�%o�����d�;��/1r���Cr��+.�Ʀ�E{��:� �9��Bw{���v��ЃR,��Z|M�6��WN��}������rk:}�z��ڼ��l����Y�������>���d��߳���5�Mj|!�@Q-P�ۡų;��5�<	-h�,K��yM8��0�@}͟� u>}�)�ME��`P���oz�-
k��:`(ix'F�߫�"""�jf��Ij"M2�B$��/��P��3�J]pC!�#���m!Mf��*g�?̍c1�\ c��!����xO�r3�.S�5��I���lRگS��.��N~F,�*��Sȷ�l�*�)��Y�l����	�L����{B��K�y��a[u=�f$�e�d�&FWt_�-�_|�X��8~Su)ㄎ�0l���B	g�����E�.\F����� C΅9������z�b�r-�RD��o��QDΥ�E��) 8E�b�J�&��69��T��~ź����KiCN��%c1G�<�F�$�ʬ_x��+v⣗\>B��z²ө�h|��� �,ƀW����3�%B/z~����]|i#U�1��)6B6`�}/�� 5����%�j�O�11$������yC����o�9�,֣Qo�hZ��@���N-�N�Jg��q� K
��:w��}b"\�9d�R錡�+߈>�R���kg��h@�|�$g�O��8M�K#J�V<��4�o'�#"�2���KFdٵ�S����L��/�ݦ>��������c�$`N��:���`�[lC�kY����Nظ�O�XMN�D��ҫn Ɣ\ܯs��A 3|]X�髎Y��,���K�&������Α9/}�'�ɭ��ʭ�Ԏ���N�`�����_�}��^/I���ƪKm�v�l�3�k�c�!�\��s�.��KЁI3�����A��2��5��vIy�Y�_�E̫�eIy?Ϥ�l�e�:�~`���b�v��Ȧ��ɵq�� �3�Uɭ�?(f��1�;���A�u�.�Mf�����Gr� s낙��smm�-t�Q����=e��S�%c�k�3���{.���������/{��=fLm��+�~1��9�2�Nc*�R�ţ��o�9� $�i,�#�rӢs����e�{��o�i��&}G�:�N;C�8�>8����G����d��c���ܿiM1-#�_I#L�&�UB��� lk���X�,t��d�D��lh	k���y]v�z�<}Ǭڛs�;CkY#\����}��gs�z=g��EM����V0�٥�Z�Kך�����.�g��x��c��^�w�q�[�*6�U]g�S�Ig���	Ȭ;C�D���?~���ml?T��9�gR���ǕX��-vQ��qU^"c4�}::��[��eɇ�D @�^���Xa�g~�
�g�����H�v�ݶ�N))���:?%��u��zdy��-QQ���`?ۻF�HC}R
=��]�����h��<*�D&wմ�U�Im�L��^'�Q!+�l���cQ���W��]�%1H�m�L�8�s�<�v��͜nk.�� ^ ��B+�-k~t*NWx�~����h��v�.�4�/a��9>UG+W��fz��F�#��˼�,�X�D��u>䜍$�o�up.��02ˠ��� ���4*�VW���k�*&M�;�_u�W��K�2j����Z�,�5Z�VKI��:��ԯ�rWCu]2h�pEs�xk�pW��4�-CyX��۴�r��`u����P�'4
Kj��I�b����`��ډ\-��U�YK+5�D�d�?'H�'�:8�.M3Jq�H���Zq�I�8�%�Ȕ��ؗ6�DӦ�W�k�Z��)c��g��Ք�$�\QΌQ|CN�cV��dZ�b�[|��sIJ;���W ���%J誌�3-��Z�Dz_3ZX�U���n4�B� ��U���`M3T�m���@��yǗ�ΰS�������¬�Ii g�30�@���9?���S�!�`}��\#J�Θ�l~U�B)A]/�3[�߿�j��bP�U0�z+���"Û��Us3��W����h9�+4�����)�*q��A�Pz�p�<p ��*$�r("������'�BѷO/�$(=����GA*�10`׸g��7�N7R���[N�V]�Z;�$277'�F	V)K&��<��_%b-���I��<�c�+qD)����~<�4h��Z/z'���/���'����C.���Q�yG�C�r��~��%)���ωP�%3i"P���!ӛ�d�����������#s�܁V�,
j��O�p��rԳ'{�q)<Ô{�rd-۾�(ֱ�y�i��H1�5
4�I�䎶X+�L*>�hue��i!^$�g���_nx�b��%:}�{��M���kO���h�0Pؘx��J4M�4���kO(n��y3�V>����=��L[]�v�j��z��H�U�Y&(�4_x��� �b�c�F�K��`Zb!�݉F&Й�l�e����|�a4��5��ajV�B�Ky]{�$ѹ����g[�Y�������x���Ӗ~�<�L��X���Zm��o�j-<��[�#;3,w�]���<�~: �v����!`,(e~�*p��R\�'��z3�>�RW7f�g+Qˋ��Q�<������6�fD�<���~\ś��%�T27�(���	.�T:A�ɞ�e*k*�Ů��Z3�TPZ����$�5�ݳ]l�gF���9~5=����V3	�ҝ�E�.� �tbR�xP�M�|��_����I��]J��r����A	�����J��Bt��^ނ��B�`j���dmm0}t��w����^A�_����q��~����sx�~w���2��q$�#�?;��� ���o�s�ƥ����H��[�/��Gp�U�x�)���H����r�>�S�4-��Nv���mE���-%�_#���5lX��~�{/������[������s�m��I��{��7�i��]�u� PK   7��X'�Sz�  m  /   images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.png�WWP�E �$�.��(U��TAz/�J�.AzI(FRT:"A@� ����P�j�b@�����>���93;g��즚�2�x@  �Y_O�좺_���"�\� ^`��m p����ma~r�ޱ	5�E�{ P(����o��K��L@���-u �対�-��|r0�����|{22SԈm�����J0��d�]��r�2�~�:>������OT��9tW���,&Z��IB)����Me�iQﭹ/��G�����vѩ�6J	{NԜ��O��:(s$|�T��a�k�W�jjn�cX��e�!|�1��/><=�Q�����uu	Z��y˜��{����Z�xc��8ЮP!�Pݏ����]��J�x�nUz��tY�KD[N/�!�n!h�t�-�)�ZT����HXQھb���3f����cn��r��:����?L����m�?����#"�_B>������+ń�N�O�	'�a�!S̡�ɳ.?�K�+糮_�1zU.D��R��s��LM>������IZ�Uy��N�ʻZ�=^1����&��/�j�{~�B�6�$.��h�	b���K�
�Nv�5<�5U:�ش��ґ��]|dӏ`U�]g9N+`��&\g#�&0Ii�~Wi��qF��G��Z�ɻ�<��=F#P��{�q �?�(/M�fś��&����ؖ@��9�C�L�r�KV�%���gV3)"�r���9���A�1��K����&�̑~G�ZS��`����z�@������2\c�)��u���fY�U���J��������t����N§��r��n�DT�ם��I�4ca{�4�R�/g^�Z΀����*�]����6��H����4�����ђchw�n��In�9�6s�kž���s�_�q*�8lJl�$�B��J�^!���g��YGTW��{�Y�Kv@�~C��N��p������:F�I$�y/���=��}e���!7	a�y_�,D!����\~��G���1K���۽��P�1�^���K��]/��gi:)/DT��ձ�W��4�e�����׻�TP���N�Ĵ�{�|�~+� ȿ��TfT��_v�]z6\4�^�(�/�?+r�^�-�R\+�d�߮��`vͫ��I����R�2���#�:���\���/����2~�ޞ�6�OT��A+��U4 �{��V�n�L�9]	&u�Ê�ʁq�c�IW7F���&�ڿ����:�}؆��٣��C�ܚԟ[k�&��>4/irƛ#r;���?��!�:�Q�n��j��p<�@B�0�?��`tty�j��~�✫~����]�͡����}�`洴z�hw�S@'2f  ��!=�7��r�\�pW�쨏����C�����xI�����TIΨ���Q
B��������������D٘!��|�^���t/v��_��M�����-9
�ںmE�m�K�
��{�(��yw��2'�y�4)K�	�WN�4{~G�"��p�^T��W��z\O�g�Җ��N��?��g�g�a6j������o{��xq�VD���r<Q�R�.Fw�����X5�͑�wQ�d�@�ݕ�0(�!`�5�6�8�.HלI96�<��X*����AoV��W_������ɼ|����.$��ڎi���J��Σ��j?��1��Ս��tƛ�|�;N1b��3c	e�~ͭ�W3ɾ9�2	4�';+�~1?מ�\np�E���@�9���4��V	b[>tҗ�Ψ�\n�O�G���B�$�ܯ��l����bH���r�(kDJ��o��������50qu%�Q&�l��q
ah��B$@��T�>3�=�KR�a|D,�'�RD�7[w��p�e�	m�`#6�-�z��/�R��I�A�S�ݥ6������H�G������׸�<Ի�}͒A��)��?iS'۹�dq�@0�p���s�uD�EJ�~=��[����\���Ű�˺U�Q�>�N=�)ߡ��h����Q�C�t�V�g4���5".TkN�l[���?`�z �"�����9�� ;41�r�0Zv��͝�9��E����hth��kK��iea�a'v�/IT����"�R�aQ�2��Z7�M�(�@�8qf<	҉x;W�+�\l����?��߫�å��^-MW��<������:�[��(�Q���h��6@�2zP]A<,��3���F��[��~��6͂�J>
өQ�Лw��z����	8��/���M�W�n�=�ѩ鮎(�O��N���'�bSK���%��C�L��M*sޞ�嚖?Js6�.Hz#�o`�]�k��Ӑ�J�}�gA������N��[��j�
���&�u�Z���,4K�:&��V����W�����w����'dӧT(��ϏvpI�1"���ԥ�[�N�C����l^!����d��[N�\�������y7�s�������!/�B�'S筱d��(
�f�Lc�� �ϕVG�֜�y����Y�W=X���C=O�x�?�}�Ͼ�T8Ab���'�r�}����+n����o�8�n���Q�8M�ubC��S-Wׇ��Y�Y�^h��K�[���y'�>0B

�U�d��� �.Eo���v�[W���
��mYe��>=Gc�ְ�36ꍽ�J=�U1eR�ѲoR5�q�DL���>.o�ps���t��&�V$�P���s��H�3s����t���kJw�Ɠ �K��YK'}4�����N�; n������`��~�Py��S>�_}�ff���{-��h�YwaPg���UAt����#�c@A�τA�5G`��{� �'an�')�,�8��&���2�>*BaW�c�C�t�5�0m�niz���M�c��I�0+�Ԭ֢7��q��H��d;�s�~��q� ������83�{�h/�#��nC��H�߳���v��M.�����l�ýM����,{�	�!b:@��LN`�gIZ�I���]�MK��͚o�/ܨu?�Sj��Wbo�	���ԠJ�1/f�S|����ۆ����VL�
��d'�ߩ�y��
��:n�P&)����fb ����T��>�W�Ŋp�/��>��R긥��O�9���W�J�W;�Nff��^8%�Ƿ��R%Ґ��&�YBi��3����a�����r{t?�)��⺜�D>��avN9��/:G�
]���i�alMzy唣���>2=v��"�DD����MG8�IYfڑ@:��?X�:��[t�<�MT��h�v#�lk�.��k��j�i79N�n-N�Չ@�ۇ��%
���!ˇ��&�M�i`,���/���;q�t�쩉�%��v���^���`5��o�½���gnΓ���W��������5������+ŗ#S�k�#�g,=(�.o��?~�8�~PdbM��z�S�Q���i�v�o�ք#���Y|�n���xSS)P��Kq�1��J0D����[Z��u`��Gmo�$}�:����8	y�;���7{�?Lg�w[��w������__��;�1A���M|��gJ$[ܣ��w��{��M��&�-VL�FB@�L������5��_/D��{9�|e��\�s�i|mx�S��9i��X�z���R��%�sہ� �1�l�]��5�^� ����ɲ�5Y9�9�M�G�V�׹�{����Yc���7i#���T�S���Ų?�D��^�ˌ{>~�!��82T�;����ਊecС��D�S���W��X��L�/PK   7��Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   7��X�+�s;  z;  /   images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngz;�ĉPNG

   IHDR   d   d   p�T   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  ;IDATx��}�dU����z�B��=��ff��a� E��~���bXu]W�[]W�.:,b �H�!ϐ����=�=�su����ι�UuU�V�ou�Ztͭ���{���p�S^i���6���-��d~���q����n�%�c)E�Q��m2i�΅��Xi2S,��'m��.�FQ���-���Tm�����b0s�;B�~����e�>'Ax���;hW��������߾Om�P�-����sC�z�C�"�"�ZȐ4]PR
��m����5�������(|��D�>u�
e�ڶi2O]�m��$��0���9@m�������+��XҰд�OP�1,�|��� ��r�:�P�����:駙9E�)�3��5Pn�H��~{����mַ_��|���O[�)�٩����~qme����
`q���eIm�ō��!-o��/@Zє��7�dڶ}�|���m�
��-��!��he��x��u��6�o��~������_�$�.Z|��/LW����yf�!������o���h}/�|s�o5$��`qQ�)^�Z�,�̲��n�V4��8Ǧ=�`���e��J4#f4���`ZNѵ�iM4�h�Ry@��Y��3XL��Ч-F�����k6���,��LW���a:U��!�����
�<�.�0�x��N詔<�Q.�f�dw@���H�t5�C?z�v�f�ॕ�g(x����sYRa��]�^��Π�)�Ѡ�fF�Y�o0��C0��+p!�h�Iv;�H�8]���՗
 ڟ��h�4#��H���A<v����A2ɫe�{��caV(�(�Qiy����X����3�W3��@X��?�EI4c��j!]�"�� ,d}�D׮[涯�xSԥ
�3�2�b.CZrbe,�2i#;}Ƞ6�d5k��x�X�F�`��h�o\i:㼹�o�K/<��4�Mc6�*�Y1�g�b�)�L��E��>y�يܺ�652�=/�P�mWHa���H� M��Z
3�3B�����h'K*Mk1\��cC(?z of���.j�X�d�X/�Y�Ҽ���n��iE���1kD�͊��u'�_Q���n8��c�n0e��ym�à]2��ߊ�T�u��=��,�~O;�;=�K�n�"V�G�VB�zR��GV��D�q�[�Y��[.-n���Y� M���1�%B��Y�R3���������Ĳ&X)��X�X)\N���8��������{~���*��X��4#��j藃B�dY֓�P�6�t�H�����f�̥��>�Į�M<�U?!���|�}˜϶ؙ��<�����6��p҂���nz(CT��>���]���߲����[�D�چD".�a�.�߇v3"�8!iU��[ݼ��4j�9����#�x귏����c�觕o,}~�1��WRʂ܈�4�m���$/Ȑ1�6�������ӏ?��J1ޱ��,�u"1":���L��qO�Ik�Ѯ�!:�PuY1��+#1T66b� �x��)�E�z��P���ebJ�p!�BMQY5�=�@_��y����s1��҃ŭ��՚-�]��}��`�Lc�4�E1�8�hV҇6{F�+aAMezN��J�Lo�$�]]���u%P3,�)�c�D&����&�������D��ٝV�J���54���[`�B��2f�V;m-k5�uz0�?.�d��8M3ᯮ��ӅvR��OΨ�l^����C�3���'�(�Hf��,�o�&�^�n�^y�;_�n5m��F<���*�d�[�8��z`��J�`_��D��;��!��VRן,s���@g��p8PQQ!��O��eg�����)Y(��;��o�.X����ΚfX��0x	����k]#�k!;w#�3�:넥PK�C�`���:�E���=S\\�?���H*�Z���Ls�K&��H�h%h]ؾ�!<���(00�L*-�|1q50	}�82� ���X�N����o~�
�;C��W��";f�A�Ě�O���P�a�>2u�R*QP�c+t{0��|r(�F����f�ʈ�g6�^3܇�ۿV[�\d)n���e������Շ�o�C~4�r��U$���i�%I�T���좉�!��:aŮ#�#��Q�%e�����E���}Q�����<�h����4GؿEE"qv�ˎ3��B �%s�%�/- �3s��lᕖ`+�f=+��i�\f����P�I�ξ6}��-v~:����-�CH�&�|���{&Q�b%�z{�EgY�:����:������m�ɫ:��x�x�w�'���]�ǡ�*�t|�܍k�����F�UR`��K<��[0����o��zW�>QgGR�����'ahC�=�ъZ����Qd"���z��ƞy	�?7	�Q2��C&6������ߠ��sz�p����.���HX�2q~>����Iv�2ы�Ƣ/�'��g��iH�;}U�V�
��t�H��)�����0r3C�0������$��̶<p)�m�o�9hi�HN0>{Y�����E��CB�i|��jH6R}'�����4A�kj�*L���V^)�(��a���O��@�k٢�$��5@'"9������D°R{=Grt �8�d��Zh�{��TYEmbЏ����*�4�3�K�ӥzV�Ok_h�� �B�A�C�n��g�gƆ�coB��Y�����j�7�L�����	�W�L�c�]O���m�.[����u��P򳏣���a)��؝�G���!����|U�y��ct��H�1$b���gP���g2��?���J�$������-����v���'�p=���^��@/��%p�{���;܏�+އT�a��䋯��Ӆ���,�u�QMe]���G����:
^�!=Ǡ���#���,�C�����X�H�UP�e�p����lM`5w�.\.�f
7N:;(�*e�I��I#�JqzR�}�t��S��B�ij�V�DM�O�����]�@�O�~S�Q�-�
_K�*�O��Y/�Eu�?�pԏ�6�c1�%��t�sa<�l)�bvH�woC�?��.+��4�.�i�ҎE�J�5��@Z���"�=��Ϡ�̷kl4�IHU.���v��t�LP^�R� �i�T����5H�hB�:!���	!XH�����-��ό�BO&��0��#6��C���T����a�R����Ӣ��	Ȓ�>Mb��!{�P��nc�)�,>3$2��i�fxኘ�0(Ғ:Ns;q��C!��yU���S�c�7����k"@3 ��4�ii3S�y�Nz�J�X��e	v�"`�;���:�B��
A0-A��;��7"��FJ��H�B%]1y�� ��Ĩ(\OO�c�G���DL��J�[�x&�M0I�F�X�'��oC���n�`�D��L���H��hZ��	�}$@D�т�1��y����|4J$#~��I%��f�"ZS��� >�>��UM����f����v�_Nm��5<��`�D�'�UX���H��~*�#�l��*����C�o<uJ!fRC��0�K�����Y���ob�F����cV��?�=�x��&��e�~��%=
3#��U^�:���ue�8�)"��9�"��b\�~9��������i����7�?D�_nw��M�L/��M��s���s��9;d�P�=�O8V-2Z�du/FN ��_/�ȱ!�0՞v��}���%Bm��ϬϨ�0�zF�N��GF7��r�i[8](�X��uE�������$�����O~�n9c7]������Ӷ#��au�浈%�L�o�Z�E�$&�7�N�Y][��HN[��� 95�W_��	��c,>�N��w�����n�yYhln�燈����k���Mm��a�/&�Y�q=�B�lFt��z�G���0�g��9�^���f��� �iaC����!۬8���9h��=p8��$@�
��h��K������o����VU��uo�R��[i)DШ��d"���
�k4{�f����@����Ց4	�z��ڲ�O�'�E@����MŨM�\�v���k�ꢬ��xt0���T�(!�p�ظ}��CH�;�g�����,����K���Yh���!�ӱ��t� �L"M%�CX�*o>�?��C�y�dt6�����ק����g����eE�>-���/������x�p$f�8����ԑ� ���Ț�!�+��	��ʜv�=Dv����N�|�KA���7�B�1)�ljNQ}�=��;d�!�H���3��=���@s$�K�feD�f�C$FL/ll��;����V�<��7#�XN2�˕v2jB�˝�@�����D��k:��߷dt=Nl�p��\�5&�tQ%{|S��3C�sP� Ms�Éd<1�������d,mY��7�wS�_�wi�w�4��~�~0������Oi�Y4L���%�00HD�&R�F;�s�"����*��;�}���e����v���'F����f�&�_}��}�:�Ēp��������n�IcwN���:�r2����l=��X�픭��２�����׊>؅�������쇢1d����1r�LzA#���(�"�P�u�[�!,���сa������rܰe�	?��r�B;�Ey��a9�t�cU�;ػހ�؎��!A#�$��meY��s�5@����2$�	bH�]2�t�1c����\=�	v�����;��=32$�}n��a��ײ��}q�"��8��
�{��@������1V��@�4'8Dk���o���",;��-ȹz�����:�A~��ާ龳�!|����v�a�/ːI٭�myF�$��bV����b��w����A1CF3Sǿ����
s�'��?%|O�Oe*?v��fq��e3����-4���F{���>���^�f�_�������2�nN&S��=��b�,1�E�����F�B��b��n�Ӥ/��a���r�v�z&^Vp2\�2�'Ơ%�0Ek���ԊL$�����Y��U�����@g�^���#�u��{��뀕���2�#ƭ,J�}Ub�����R�B�׳�a��HRȯ��"���J���$�����
C_�sti��2-9$�)��UX��k��D��vH�D�}��C�"r
e�\���F�H�����.F���_q5��
��m@��qq��K�@���&�x2g��E��h�_��I�\04W)�Vݢ��(�{(�� �~qY��y�~�5(�{ 0=��`��P���pd4��ë��ِrb�x�LJ��W�vHn��gZ���Đ�e5,En��ȁ��\�$¿���h�I�7�#nm?�e�����]t����!�~z?�'3��hVL��(+�'�'�![&�Q�����PgL�f��~��AKP�@.f�Ёي6[��\�~Y��� ��K��ٞ"�'q�z����Bv:Qt�F���?���W��l%2�\3�r*��������)l�횋��&
�b�|6��٢������I�e2��8�W�2)5�XA.dk�������0���,>�\�[�b�W�@:�l�Ӫ�8�!C�.��]P|%P#!�D0�³(�~�����
{0�QKƌQҴI_�@xYhN4�0��� �(%�BɆ�z��"Y��j\ͫ���#��+p4��:�t��u#?���V��?�A��v��(m���b���#(��5��p��'VW��?$¶��8����Dp��g!�櫰U׊	ȓ�VY%Dw��A�ܙ0� ����m�VQE�"7��ar��L�@WS�@FB�Zb$$Y�s��1A�Ǎ�l�8w޿�E37N�1	 �z�D���C��XfxXYXD�XQ��fأ��Ӌ������G&M���`	b�ٽ��	�[��i'��:Խ�dB�GM��ޤ6g	z�{�i��썶��iO�<t@(��Ѐ�<�N#������V�
���;���$���[X:�z�ɈP��(�w͜La1�Ngo#�#@���pVz�a�Y��ٵ���2�cN�هk7��F��wb����U����H��B+�1�� �1%�oG���D�o�V��.�/��s�a�0_�
�e���3�Z����d��ayE3"yi�y�V��AݎǬn4�^��[����E�"�cq?~/��2:;;c�_V���w�Ia��~<m��Q|݇�#�X>�vZ��|�k_�/cC��=�1�G�B7�T,��A��r(ⓗ�gl�ǯ�n�:&,Di#��L�W�G�n���?�{�)���"Z �a�i��amA����Ah4I���'�4��p䅃�R�(�P,L�J�*�|�g�A<V�̄��-�i),�憢-`e��f������^�+.�^"\6��g������><�������L�1�q��V=����i��W�{��N�����&Y]L���$2v��D�B����C��'�Z�] ��
;Rezv�W��-H?|nR��6!nu�%{�T8��=�뗠{Z!�H@=F��ƿ��+�<�V5��	�3*I�S<�[u��ۧ݊+;����DҒ�2�� �ǘ�@~G1�~��P�?���9Kt8S1�w���x�[��~��⋌|�drF[�ۍ�r����b�)fw	�X�f�Kb,��C���aܶE��c/l�r��c>�b����!��C�¦�{�|��HZ�yb��V��p�57N#}L+��9,��}R'��>$��ܷ�����k�M������ʍh��M��'0�ė���-���3O}�8�u�pa8�"1�����%m�`.�p=3���'oڄ"~�9h�h�ӆ�n���>M�L�q�	����$��_R!]��5lw([�>4��<#'�K���6v�JvY�hʆ��
��꩘^6��>J����U��'�)�$%Oޓ"�y�Wx`�bC�V��eZ9�2��-�W^u��\�(Y@��сM��b�E��х�9�f��!M�C����ڇ����a�V�qZ���c�A8�[HIy��@�	B�_�S^J�,C3K�Y�E+��bS eǓm/f�*$�����6��d;_l�r] y!��?!�0����g�M��9�4pk;w ��DG�+~���tE#}�o��+j��	�� �(p�%^C�=.�Sߘ<�@�Y7Ŕߡh�W�ؐ���%
B_��͹�"[�Ղ��}E4�{C|���p�Q�dВ1X\ޜ��=�(j�:�&�XYY)`��~���	/��"�2CfIr���`E� ���F��w���;9����p(�7P7N��,%���ɺ��pVT�}�K-�U�\�>��Ŝ���0;6	�{��%dx}��_b�m/�ɑc�����,8�>I�e���R#1����*w�\(++CMu�	j��̙���ƻW�p�d�$�h�����'�R(�x�ڍ� a�A�rF����ņ���`�ß�{��<�JL�~�= _x"0�
N"�ԣ�#_DQ8���/��D�\9�+#!�]�E�2��.��d���
��p8��H���c�/ Or�I[,EQ���x�C�#�#�%��=�Xk��bt�0c������5t�n�v䈱`��K0U��g&̸'��tc�3��D��|����(��:Ay$�e��хzlJ+�EO���a�H�����pCQ,S[60�i@D�0Y�G��!f��8󯺺5U����#����h����Ç�q��֬�v1��*2��xb���21&���o3�~�, ���֞��}�8�2+�زb/J<L�4<<Hv��N��*n�?X��"�,p��!UUU���LQ$=I�B]�BkɴL�k�	��-R'(��D"�λ�����+�PRչ���l�%.�,���B3���hoG�"C�|[+�o-��V�sX���&e0���{:�%��԰̜?3z�V�ɑQ\�e+"�Q2��ˮ�h_m�ˠ0[U#G��{��̲"]ŵ��7^Ƿ�������[��pS�EL���FaUk�1����ۈ��|I@� [�Ծ��ń�M���[n)@YYg�0������,1��Ċ�8ғC`��۲
�S����E:�B�Dn'��GM3�FY4.�ˍ�d���Uը��Ĭ8���	�&�U���f��b�J7?���d�󷏡`7\֮]+c�I����}xf�s(&��,�l��l�㍞�4�5��e���@g�S"��}Y�#X��0���(��*����`���;	�T��d.I��4��@� ��P��]������8����F�57>�������>E�8�����Lx���!�Z�
M�a=�H�����µRc�#u�PS4�Uh�i-z������/��T���F��~�`��b�ϋ4d`` c��|�=Z׬1|\s0�Y�q�Dx�wX-� A���7�N�I���	T�!�h&O�m��+�*��[s)uj;��Иe�p�Y%%�������8�����~�H@�0S��q>��=�^{F��`k��\B bU�z�n����@U]����
l�Q�����"�W*.���D�*u����&h��D�z���3W��4F:�	x�⢘|ԟe�n����*�X%iى�{�xz8G�*HӺ��j�n���2�/L�"�Yb���8�&�M/̈��^�S�I[�I���ҁ�"SXI��e�S3F:�}�#���	|M9M�O{��]��4S�؞K�еե��|~���9��4�	�zpa�	����:��'�Q�NzM���l������.f�[IR�$�.�����!�zc^��Z�
Ȭ��ŃH��%f�[Ҁ6��Z"^��Ļ�}�S�np�EƲL7��PL6�H&�Ԝn�̭��s��%9����"�W"�����>�n�B�m�&l�&��<Y%�c��/��ƅ$}�<76���ǡ�3��7�� �Ua�I�����~�N6��[�R��a�<�^	��):�O��}8j+B�KAM���(F�:�*m9^�n'n�����p�ھ����Ӄ&E���2�W#zp�'���ߋ��h��ۍ`�	|��# ?��ag�x��Fr'!\'G�n>�p�x��L�-
��FFFP�~-���j�oWz!�IhW0~��aTUV���6��MU��?���M�Aó����7X�В��t�3���>�I��`�-��a��j���c�h.;����a�:Y��e�Wxx?�������=d�0�a8���|�)A�އ{t'A͙��YtG��Q�i"
;;N��|@A�P&��:E�IG�<St�2��|4>��b:A�k@(�0��DC��**��r/!}�z��ć�,Q����O�O���&K}�=��1?�)��p�s������y�#�8A+㹗;e�w;Ĕ���G04�4 Y͹]�*xq��Z��>.ғ\�Z=|P�K�rx9��l�_ºj%��<���ݹ�!|E�D���"��Jp�����&{g��{��9��� w[{��}��dk:�O�'��
�A���A�P19�uB��đ+pP��JJJP[[+���ȉ�jG�E6�<��|���R���&�1*�d����OJ�.H�z�
]$�͟��̨&��!�:Ja8hL~�����;}�L~?�L��3�!��8qa�'w�Y6��#�����_Ax�F��4�������L4�e�턪&V��k��N����Alڸ�_v�ܱ�>�(���66`���@��.�9b�X}%�^?��W�QRQm�(
�$<�.!㩟�ub�h*���j�e���+���#�����\e�����E"�|�>LsJ�M�c/��.,��`I���C�xP�_�au"�X<dHB3�Kl#�"�;���՝��34�Pz9M�Ёɭ�D��Kn�-[�o����.l�$�b����[�ك�^Z���G��P�����=�z��`��M��T�JZ����N$o5:6�[O���}b_���+Ѵ��h�x�U�2����=e;��,�d�`Ög���[C��~�$I݆h �FZ�	}3y�\YfH�~��L��$N�<�#�w=�����Σ����w�p�͂<�椩�oooǦ�N��%�}��b�5]�ޯ�iSv�p=�ů�g�^{�G��}�qU�r,�4�e�d6C��T��6�uB������'D���&�E6���14�M�P�#�1��*���g����fiqĐ�-�səL�����	#���iF�S6�['tF2�p9{���c�Qݼr�V���C���x&����g�_��ݮ���\�"T3��=b�o�8˫q4���چP,�DA�a�l4�W+	\alR��#d9��������:>t@���"�Y٧zc7���jY���Qw�����8����w
Ĕ�;Q���Rz�%����V��N�(Ny��{�J�uv��!v�gl�"�w2��+?���"�/kF�nZF��>�Bg��\�ؽ�m'��ϻ�x�`�F����� j�����
�9=ة{jjs��J7-�GFe@1^8A-i�1x_��&�1-��3�5�l=KlSQL>�4<��F�����M$F,(jY�T_����G2)n�8�H��@O���#�ۀ�@|g���+ϋ�
����!nK�Y&E޸|�����>�gt����Ҟ�獻�%��J��)���g���:Z��Hϓ�i#��X��o�.i�Wu<��,������蓄�톯_2��L���[$sv�M:jz*0�\�;׵""�<>��\,E�[o�,� C=��C����aD��`�!��@"��BǏ�H�y"P7���u?�G��pM ��S�˼�e���Fq�v.Ab�cɮ.���n#��!+���6\�!�^���$&�T1ƤQ�;t�C��=C4=��+���QxRQaq�R�s���=�:'iZ���[�l�d섽�A������u(�����dMK��J2�q�1b^�9����Ȟ�#�W����Қ�:q�
�q��%��O$MM�ά��i���x� ���	z�]n��WP�U���v$����b��P �w���%w<�˗§�IZ(�+T.ݶ��v}��O��b��^MR"J�]�+क�	؊��4{ݰON�E2:v�؎�&��(�B�f�N�׹�T�[OB���H���-kB�d��\�lTo1ĥ��2MԨ��1�Mے͓���0c�o~9p� .��,�P�n$��;O822��=>�.���J�:W�3!r`/�$�#���ZS�T$*�a:[�����!��4�Oı1��/�U�\���~��.x��Ι����v�vثV������?*�Qݼ =|5�����q�kP^���ŞF5F�՗s�#���{ϫ�QG��b�J�J��-^�3���J������*D{���E��R\����)	fV<����N������b�����"$߽[����w�}~�[σ�3���?������>�?R҄�n����)���	f����[�
S,���'1�%��r��r��mr�K<��r�6�S�y���c� 4;$�8X�<��� 0&i���?Ɨ��c��|���ouu��F�ܫp��X�Q���h"�,��+���z߻Cl�)�~´J�6��!!N����9
�(Ь����8c����/�燂�V��Õ��V�E�
����bqó�\A\�j���&�����w�,2��kk���l����ϣ%�%`�d��0�����!>�����y��D'�����w���s��>���p:��M����[��Zojj��3�YGɱ�����[k)�+�ov����Q>6������4����غ��<��X���-JHS'�H����Ŝ5<uޡ.�ϲ`�D;���`ǵ�@��Ni������POn�c~"C�H�ߣ-�{xX�>��?���ċ�}%#����
��8V�g�Y��8�ÿƱ�n|���ओNY�<Ax�d0�ǟ~/��Cv�W�ܣ͒�Ęs��/}5�ӳ;�����5��[��}��nNv��F'o��ྀ̽s�y���H�Q�;=����[}����H)(���o5�!��J��H�1�ɨ�Bh���0"�Bm_%��co�����W�2
�3�g����뱬��'wubt2A"vj�q���"S�"�p������GCC�4�]�������H�h�T%��&5Ǵ�[�DL�N�\V��V��kO�ˌC�/��T��N�J.��.��|1���nCI篰�p�8�)CW���KkE�n!���`�-��Ѩ084�~���wC�"]B�L���g�j��z�2�#�ܗ)ű�w@"�u*�0���7� ����2�f��ĔS��X�j� ��{L��s-湓�D4��]9�jxz�{F0H�т$=��컛&�
p{��Đ�׈�-�rbf�<x�o�ג�'S�֪
�%xxx�ؕ~୅�>H@`�.>���"�S���Hv���a��˅b�/3؉u��u�p�}⁹�����ԥ��V��Hb�}�rk������$#AB���1O5�����n!)Kbq��xN^�Yc0_�����Z*�X���l�t��!��.���^ ����rb�˛��ݐV4s���,^���&^��o=.H�{HR�y�Z��� ���9�u�J7�у��Z�hʐ��م�"ZeV���4�d`n�Ԍ5��3b�F��S��S�� ��E*?G���P������˦��=4�Q�ԧ�:D�w������01/.[�=0:�	������II�e����i!>�ה���5��$�1E3�2��դ�V\',vf}=��+�C]���!5��!J��o����^%^��o�.|}7�)%�'�@�h:�}�=��P�~9;��_A��ԋ[x�X"�X�J�����I!9����O[����@H��,����Ѹ�L$11a����,����pd҄G��IBN���"@F*G�,�XWg�{(,��܌6�y�t���Z-	�$�+��_�u]����Q��J�af�n�b�rb����Kj���̯�f��9V�"� ����@?�À֚��Nf$�)��03Z�u���{8���&ie�=D��_��H�S��Ey�6fF���A��/6�#qw�/g������z���p�l�ĺ�:���rPkYC�@asÝ�Ƥd�hξ`�7CK���O����<j�A2��Vd72�x�&o���k˪�%h�U�S���4.�[`#��&�z��T���*¦�H�z��[@c�j<.�pXr�}�b,	��������mB)zV��.�D��{Ǆ(.�C%=8��Wn9y-�����`Z�����eZ���gosh��R�MZ��!ۀ7�Z��;�$⪞J䗳kO�f����]QPJ��C𰴴T���WI��'�$���Cq+�	11øp�>��9�<���J�-ƓP]�VA�ׂ��W�U�}N�Q'�l�h�NXeS.��"��yC�@Y�?ہq\��f?�z������ET1�.o;k1Ђ�>CY5Ը�W�;V�-�O�<F�W�31�ҿh�2����}�����w��V��Ob��^�$��I7�����Dk��ܲn��د�DVn��n���K8W�&���w�Wހ�<⽯55�Ѽn\�R�߭��O+���B(k��k���r�D�-����)B5Y���G�[i���z�O߄3�p1ڡ����E�YMm%�VTQ8b����X�B*�� ;����I����,�Be^�'z�i����l����al�#��<�.흃�b����q����
�r(�t2t�3���Ca%[G�ض}ݍ��
.!yG�u=#�]����~X)��l��.o�U׊�B�3��S�.e�H�Npr��A��$�O�/Oo�K���P���	G���=�����xd2��[��U)A����C�2��e\���À3������$z��X�:q��d�P^b��t� ��G�f���V"�d��#�ә�+ԔP�)o����K���7�k�"�A��~�zACS���$ho�3�q���.~��KjX~/M��km�E�pޣwuؤ��c�W�V\0u��� ��IؿV>��V��SCp�+��2ـ�᰺G���BmGt�V���ŧ�,��&nk/rQۍh?8�J��S8�����ʋ�9m�� ���D�~"�l��E�E,�~R�c�e�H�ץ�Շ,�ʺ<4B�.#��M��&ɻI�3����Z���v�b�b�c$	4e�eR���5��}�m���~6Ĕ���^�i_���O��Ж��fb�&7y����c�g��$z�Ľ�ޏz��`����#�ȐcCLl�5N���ࣻ����bbV1��Lz��ڲ@R��3�1s[��m9�C�k+e?Sǜۈp�OL"�A"vS��2u�ܘ�D:� ���|.$��䤱?�&�B�L��mMNX/6��2F��ߊ����@5ι/���Ǡ�qz�S`9S�C D;FS���z��&fӜi?��|�-��?�
��m.BUg�h��AB�˃=�q�]x�tG��T�����q�\�I���e��c�i�xz�lgP��|���ݫ������� ��D��s�F��>z�7��Czl����`�&N8�','g�6�"�2��wb��;�hX.z��2V�|H��������>�H�A�h��]$����cF!CL�0��G��,Ѝ��^`�Wel�w?�'N�	[f�s�0C�$�rK�� D@�|Z�i7�9��8�ϫH)�%��a����A"f���B�4r��"��Ldm�=��OT�zf�qĬ,c���}�"�ħ��~3�x�
A�,����Z�U9���.��b?��SH�E<�h���"\��8�%���.�i$#p�*�"��
�E�!�sz�ԣ��	�=���d1QO�W��#�uςl�S�=��Y<�.D2���ȰnO{a�t͖���o�-\b�    IEND�B`�PK   7��XJ)@i	  F     jsons/user_defined.json�[o��ǿ���j��_��Dɩ;p|����\:BmQ�$�A���%i��A��H�f�3�,w�i���vӓ�n㺿j�,W��Φw��,ە?�\��fW��n�'���������]v��[m�n�ϫ��]��G���,�og�e��6XTXJ�T]׈C�UZ ��Ns[�s��u�r����P�l��d��ܗq-ܦ���8��}���gV�KN��"^�
�uE���Z�)kQ�W��w˪]�?RM�JKdD-g�![�Ij��j��?����e�}��������;珮���U�NO>MW���r�����7~.���S!�?�롋�C��B
��H'~�Z����Z��o�����Oh7�������\*�IR(͈�Ǹ���wm��0w7�t���n;�<��I@gr��7�o�׫:��^������~~;L������MN�]�v�v9���~��=F�1r��{��_���-W�䕻�*$�!�_-�����ڛ��1�]ޏd�kn?j��s��%�j�E��	1���)0^�4D9z�)��&��RȺ�Gk�Uyz���'��JN�]wr�fO�qZ�X�Qrx�&��`������/�2�����ǆ�E{�����$��X	²+����@Pq�d���A���I��槡*��a���,	�!���s�d������$��[8,��45Ea�?O)	Ea�?�ih�'
��HCC=QX��e
��b���PP���:ŀ�o��PP�iE�PR�$�)j�ß�EEc���VUŀ iY�PV� ��u5� �{�J��y�2��5���O�,�itDc�&��ş�@�(�A���e������?^��g�9"<������1/��ӂa��f�h�G�AG2�������}�E�T9dr�#GrX8���H��ɡ")T6<O�ԒPՈ<9RPB#��HY	Պʒyd������ȢM�&O���$�LpY�	(��ё���2䑅���:����s�9��v�[��P�ø�����3@j���ا)�SS+"5hO��[:[�H�S���L"R��T	�ɧ7"R��T��w"R~�T���p�<{�P3ފ����،�"�ݿfX���"�急 l�a2!/�__���L� ��.�	���X�e2�0�M�L&$F ��%4F "��%DF *��%TH���2�?�d���
�
�Ր
%6P!Y!��U��*$+��N�P`��O�T���
�
�(*��@�d���Buq�
w�������W���
�%��
�%��
i���@Y!�2�P(+�]�e���tBc���v�N��2.K�� ;՟:�6���t5�W߮W�Ý����� r��v:n#�k?������/����fY޸/�u��n0=���W��hW��V�]�oM��͏`��-ae�A��q[d��"�k�jZkf�4��!�>�p���mY~���lw�n�n�a�}7���L��we����� oֶ�W�[e� 8��rCZ�
��T7�F����f�;	�@T�,���i駣*)�p���bSS�5���uf��><��{LT����b׿�|��,�J/�����h�!UA4�f&=�z�ޣ�� }Ly]�?E�1L���X{�[=��J^�}M
1��1��C�Y[��P��QaG�vT�QaG�vT�QaG��/��}6Y<������p�ߪ�|�]�YM��UV*���֏�Ԉ˦����_sXSV��V�F؋q�`T�#�yS[��4��Ly)�FH�g�qdi� ������4%@�D�,�J�z�P%��K��LrVplȞ~��?.���ojh�	��3�I�	^P���������{+�����q�� �r
�g������]�P�a=�RɂlČVŇ��=��~���jAj\`M���=��5�_�_��6>�TJ�� q������^��:��hH�{C|h�:?�-���D4�bF)������A]�F�>��A]��0��'���A�����C:�	�J��ӳ�<EZ|Ƚv���$E:}�hA�,d��c?���:�B��>�������,�����%����E[��ǩ��(Z"ڄh_=O�����B����u�!�NژƇ�HԲVDTZ���J��q���?R;hE�K��C�C��AM�Q)�_eȦ¬���@q�p�pb���������;��R�B!j�}��_H���:���{�*t�&߾[,�u�oKGN��Y#ɉ�k��"+�A%�ԑR���wM#�w��clc�[�w���� PK   7��X�����  �%            ��    cirkitFile.jsonPK   7��Xs!��}  {�  /           ���  images/330d02b8-4530-4fd4-b6ae-26fc03cafecf.pngPK   7��X�ة� � /           ���  images/3c114b42-368a-4c2c-bdc1-509aa8451bd5.pngPK   7��X����(w  +�  /           ���� images/42266fcd-641e-4cfa-a619-b442e1b7bf10.pngPK   7��X+���  D�  /           ��p* images/5cebb09a-e86f-4cb2-800e-22da09d26481.pngPK   7��X��/F��  ��  /           ���� images/7fff522b-95d5-4303-ab4b-62aae53cf766.pngPK   7��X�IM��  � /           ���� images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK   7��X`$} [ /           ���� images/a8bb870d-02b9-45f0-bd60-404fdaa8f6ff.pngPK   7��X'�Sz�  m  /           ��e
 images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.pngPK   7��Xp>r�  �  /           ���*
 images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK   7��X�+�s;  z;  /           ���H
 images/f3037bb0-f56a-43e4-a2ff-17056f7c669b.pngPK   7��XJ)@i	  F             ����
 jsons/user_defined.jsonPK      $  �
   